��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚�rYiZ��}5�B�
u�'k�Iv��_�lE�e�C�@޹'_��;�=4�2�/�q[��9kC�}��u��HG��V�NS�?�f������w��\�q�"`҈Nd��r���F=��7-ʮ������VY� �D�+��˶U%-{�u����h>!��F�5���:!�L�k]r�Z�GZ��k������y�>mKѝ�)uul3D+9J�d��zIf&|�-�t�.0�Q`�he��ۺ��+�+H$ʋ��oƣ��2�YKQ#��1X��IVΟ�P�y>�.�x��j�,x!��n1ˬ�[iu_o�kxDD~xsqoV��E����G�nx�Z�@Ӂ(��Ǟ(��s��������]���I���k�6?Y}<�o��1a���sb��W��s��i����b��,��g �KA�j\p�����ybc���?9�]4<P�$���ZWD�HWG����kql$���;)P�\h��x���S��&�J��3"��a�8n^���tj+�{���X46�R��o�c-o\iQ_Ţ�x����.��b���dT�@��(*k��fɻNސ3Z�<�h)N���@�Jh(�����P��Et�h�,4������(;��rp-Wo��9�_:-A���R��?Ħ�a
 3[���*eR*�/D7���t��.F�&�~��(����7�А� F6��H$�|J����gƈ�b*��
�u���D���O��WYb����L�WG�4A?�a��A�M���G)��x^�9�8��vK>������n�o�� ��`5M��S>�B�M����qI��?Mp�Jn�X�K���V��k��-V>��|�3����F���8��(U��	��F1>�a&�T9��**$�p�o�>D-Z���%]L���-U[�x�S]r��?α��Z*Q����㓫�K��s����E%̦�S��!�1-vH_�
��o������Iש��%�($�,{N�9v����)g�2r72�&Ɵ�-��󐿩f*9��pL#Lڨ	L_u<^�JMqu�����i�9b�(��J�>�?(;�,�K���J�9c�-���.y����PA�y`���	b|?�]1������"t���Ҽ����SLr��(������uR$O��ق�1���|m��	�ȵ;(��A��'�e3^�8�9�]d��M�8{�̮�uFL�����.3R��pOjY��-�5j�n}͉����f�nF&ꔴ?��������.So��k�����s�Y�=ξ���'���c�I 8�i��!��U�����e��x'R����3p�ZF����nN�.��zM��˂����������F7ߴW`+,2�bO�j r`��R4��{�2�O�UF��<��޵����O�s"Q�拥	�y���S�)�©1L�v�"���uE�ݳZX��j/���.�Y0��`s�l�+�P��B�?4��aw��W�ξrȃ�'���s5Q�|�&|᠚����|�Z$8_v��ؓ�Œ�gbc&�q�]YjC�3��6��F������B�����ӝI��G�~�ع���u Ua��z��V��(��Ff�w�S
@���8��5L�6^�\�D��q���C5��֔TЪ� ��o������ad�s��l��}�
bΞb�n��.P��.Jl�1<d��+�ݫ:�8�'	��y-v��b��Z�����c�J܃ic5o��pL�y��6צ�J��)���o3g$�zE`HТs���̖�L�e���}�.�x k��/;>���A�[֡ƻ�++B�t�Ԉ'�!݇2@�/��I_�eFd�B��-)f���4�l+j�G ]��cL��*�	����t��'��d*�0	�S$����p&s�,�#3��]�wݺW��9縭@`�,�FާcN!.��L�ߑ�ӻ�UA���z{�� `����&?�h� N����KΨTa�����ǌ�R��\�u�u����v������n�;?�g~��)�O��<�̗֩z>}95��h_�K���{>�F���z��C�8� O@&�)��`6��z��Z�]fk=H.�T�7��05�'ڍ\?gzҐ���4�*���q6|`6Q<ZV)A�Y��L�Я�JFa����b�g�YZ���ף\�J��]��������O���ރ{�x��YG �G�nL+A�a�+ԂԻ�7��'�pҬ������&�
7�I�l9o��U	�w�l��d5�%/��ʚ�����Ѧ�S4ѻ2|Ҡ� /)ؤ1���nE�=�~�T�W=jCF�����[a��ن�U x��R(WeT	ם7��UG@�U͝�Uf�u��4����t�(K�?�ƻ�H�ӻJ�=j��#z-쓎�b�J]�ʂ����D�ҧs{���m���u����Jm�����zKi�9�\�e)�y�`���N#+���+|�H�F|������%-
������YB�r�{J�y 
��Q%�G�S��P�3�� �P���єE䯖�1�2��#�ہF��U-��P|��s��K���>�)P�-��esov�|�Ll^#���&�K1K:�ވߥ/h�BA����npv.�[�0y�-mZj$���n� 4�pY"/�lG��;I�[.L�y�R��WSr��|DDj�8^���d��(D��M\I���I��E^�,�R�h�YY>�%��N�٢6�&n�F%|�_x����ty��1�,B��7.�	J��G�H]�1��ƨˆ�E�M����ܓ��F���X�*{�e|�p���Ң�B��hi�ԏ3i��+��G�?h ��� ���A���S��G���͈n�s��	>���C}_�}����0��6�Q��|�E�O&qJ���[}�Z��@[������UU	����������S�Zxx�[�8�?wS���ce�YP�u�cX}5�t���WFAs��kY����}�k[� �F5�+^fg��pf��`�!�f�[��s�(������}�!�(ѩ�8�ݱ�3�E�Hn��;�x���lљ:�ܰ�Z����
�G3��#��у/����d�kt �qu�_k:}�ƥ��s8s��jY^P��tO�[gq��K�pk����(!��MZ�xڐ0 9��I�H�[cS��)�*���J��[�k�B�5��]Ib�?������1��ㄩ�pzSqc���G 5��^�8����ʡ\�XZ�ёC��Q�Ⱥؠ��_����z$�V��o�C��+�fb��
!5C�'mRɍBr� >˪Jf!j���]ݓM�{T�0c�&�X�OQd��Dl���Ԉ��An���.��I����q�oLAW��g�[e�(2u>j�|v;[Xmo��x�.�A���v�C�B1>T/��iƑ��������r�o�t�����1�M}n#��,��jD�m|h����c)yԝt�l_��%$�P�)[n�Gm��1֋n�Ca�-��L�^ѫ������EV������)�y8�3��!�m�/M�9	��Lx_�8���1���yؖl�@G��&���s�q��Gl4n%	8j|�"6tQ�`���ɇq��Cw�7���9��Ч2�r6�7z\�{��1�N��ٰب����5w?l��M0ƆE��Ƙz�V W��]����7��gi��+���o@_�~tb��58܆���򢿿�b�`x�� �&��4�U2�)\�SN��RۘĠ ��c�>�L�	��.��7|�ѱ�j�Kӓ�C���9D-yX<q!����R� ��7�:�"��#��u��*�+��&m�Nѝ���@Bu�do�b����]E��CrS�b���ֱp�F��i����殘��������k�ʨ<mɘ�����`x�� ��a��W<��s�-�j�^l�X�	�qu���uVz���qN���N�)q�XY���(�ǉ��)]�� R��pVD"��v��]����R�C�4�xA�ʘ2^ U�.��5�k��I?��@�\�f�6�A,$�q7����|�LWb��8���B�*ĦS��ٳ��`��rɚ�L@Re���-���{T���ZGz��Ԏi�W!�波lO�U�i�ۊ7-H7D0�{���ņ ) !#w}��	~�� Ц�)E��ݡ�M��@!�^���]���d��|�.�a�k����yq��(K.Y���!��FͰ�a�X;�s��8�Z�#A_%�bs_0�WG�R�;&�l%v�"߮��`;�O�֒����z�0O�M	�z�|�eu�J-m�Q�5����́��	�n� �*.�u�Zk?�d�����]��*y��s��e)�e�9�W��b��	��*��+�/�Dޒr�a�1g����ؐ*.'~��tAz���#,F��T;{�qioj	���?�}�/�㿏C������pẩ�u$�d���!l�����CѼC���0CT��U���������ݼ:8�ň�]�g�K����5�?5��0�/�Xv_���rv!�������/�+���Wߞ9�Ȉ�w�Y��=8)p����|tǪ�Q`��,V��i8%m"r�(�8���p5P�aC��H�m.B(GQ�سsP������w�2�ZA�tEK�h	c�͊��ѠTf�p5�8>U��_)'%DG�W�_��n�:� ��J�t�K^+^��k,Z������,�i�h|� ����|q�������=���x�)_G�-
����ڤ^�}"��V)�<Q;�lEGpZa��n�/��@Ap�� Wm�v��.�f�c��FM�Z� �@���n����]��z�"������i+����fì[���>a԰]������f{��y^�Ɛ��7���%2A�����o9j��)��yYo��m���� V��H�Pt�ě�Q���y<e�d�ʣ׾��u�����[��U�=��U٢��+��e�<2��.�����|�+�qo'�\��R��!`�B�!�p�UR<�:���J�/�G�X�̖:?�6�'x�`�NEc�e��V�T�<��z���֦7o>댟:����a��4A�|��Yyο�g4g����SN�n�:��2�9?�1yVY�Q�dJ�>@0Qp�����Ϯl:�3��O:�n����������1�~����:��(��Vp���I�F�%����3�FC0Lΐt�h����_�E�� 0���p~���ِ�s˭r�n
o�IWq-����C[���^�n��-ex��4>_�Ӭ�����(��M�)���~�c m�*d4u��ϻQ�wV��m�(�(m��D.Ëŉ���:P���i`,t4r��P�+�-h��^ w��	�t��]�L	�Q��	���i~�̩C�u�0Q�m���If
9����e�rmV;�{��9{������taA
2�&'^h_���-j ���ձa-Y7!���%��2&����R������J����at�홗���v��`�`�3^�Z��0'���4�Er٨'W
g}�:�VC��l��Q��%���~,�����K|�{�����@TX }������&�y��4P�%����-�����NƜf���d���A*Kpx��{�����>sIkR���+��?���LV���7*&BRjOC=��D�%�&m7ﳝeD���W�?*�>9 �, �Ґ]��le>k^Mcڳ��p��O�M���Q/�#7�Wku+�W�q�g^��!�<��V���~z�F��'� �E�=���!�?�9G�>1>hL�R��9Gߩ��l��Y�4@��1��V6����0��n��� ����v�}�6e���d�r �`�
�y�5uP�Ա�-?�6�/5D��
da7&ʲ��l��V�c���&�%;�$�Fٛl���ܣD�sc)�`���O��u�y��{B��`
����q��]/���5��w��J>vC���0e�D�q��̕i��2���1�-�M�?{���,��6�Ȍ[9Tv~D}��MFIqw�;{RZ �A��(B-���(�WX^�� kΔu����s
tQ�����I�yܯ�8]0K]	���+Ԉ=�P�3Z���AG��0���x�hDI��4>�F�Z�u#,t���$*�6��. ��9��a��AwQ�b�6rg୭H*��:���[ztB��m �c��	r�>��oC�z�A��&,2�6���p#m��#�b溝B��Nn�i|6�2���0[�uw�����+��װ�&>�б��5�́T��rI��p@r@�Ld7,/q��9ݦ�π��]y5���z=Nxx�%^�J ��!�l���&�ܜi7e�O�C��A����<�%�HޒT���@��P �+��{��%v������=� ��Q.���V�`94l��IN�{Wg�SE��ۈ0_��2-��i���7���ɝ��L���޻��J�0 V�C��}n���v�&bW�c4��cDM������L�(�Y�u�Ȁ��m���k+c��}�kԃ<ݘ�Db��y���E�Igr�X���(����l8sO[P����[�D���@��	�S�5�٩3NX�}��<��vf�3�b�Eǆ8�S~�2hF]��Y�6�pO惇����������,�8y�4� �Cll�?O���u��Ք1�lH�I<Տ.�)��!K�HdR- ɕ�u5 �v.�������}�����Ab�dE^R�dtP�
?��K^2�����w��HK��ئS��Q����	�|���^m�M;Dc�'+OKH�yT9R�ж-��UF?�{A>_�Vk�₎��avZF��^"3c����wu4#��v
��W�}<<��D�����K"A,4�8�۰���6TP|RP�O�֒)1R���gp��A�Ty�>�}����'��ګB�\���I�8�L6^�V-� xn�Qhf� �I.�B�ի�-�<�P�O��e��R��'9�Z�1�Hn�u�E:���6�c`�9ρ8nq�6!{j+���ʗ$E�ę��x<q��qo���W?i�%̾2���v�O�}����W�k�y�F�c����|+e� &� "��B�Y9��#&O��0�Kˊ;B�\�5�%.EPѺ��6��}�0�O�f ��>6h'Û��q�$E���Ȃ�"�����ώO�@\)�Z���)Nӯ8^���H"��I �f3���~����_���K/I]#-a���>�Z��?>�C��_(���7��X%�X�_� z`i+�ɔ�:�⮃Pſn��}�|j�Y]��[�����E���-��F=�Ʒ
�����Γ��P����?�QP{?�pLQI8=ļDfzQ�BαQ�^�������=�ϸ��QӮ>�I��%Vv�������5-sE���#@-�G5� ���.����"�m�Ӂ�c'�.}? 1e�s2�9ԒZ��K�$�(/��L�ߧ�.�rZ�W?�UǢsp��U�}�Ѫ��@Qi��b�.�9�Z����ȫ*�H;!4P���T�_.]k�j ��q�Y�WG�^�Up"�ĥ��9p�Sͮ��O�؟������Ds�Iqv
��5�ڽ�X;(P�Ċ���H��Ev��J�M$Hx�8 �����
<Es�W���>2S�ب�D^zX&m7ka�#�;L`0��SB�
��\t�w�qe|����B�O�鵕���L��צR��t��RwfI:����b����j����%�D����w����[7]P+��Xe���`$�������sHת]����t	���$����U}�[�l<�r�C鈰\��N��d 0߾.Bqom!���"�3来��I���u@�./t���ҫ�� =f%*�U�c�rz�o.�ޜ���͂� 1����
��i�C?�<���>RRu���~,�6e[���	��~)��Q����"D����$�������t_M;����3Q>�m(RYA�W���R�$�	��g.�����Yqj�>!?�9xm����π,<)�X�dBD�"�ߒ�j�B���me Do�_��uW�pW�ú<�.�"V�%"\"�C�1~|�@�k��B�
�ե�������!_b��em��ci��G�_�ܩnn�ntfqö%���W~���fy^z�U�f��?�������@���?�rHrwI�h���!�q���49� �W��:,�Õ���s�IF�e�)���#I M��<n/����!��s�;�*pT��}�\?D�c�Q�E�K�#����٤��TT����{�#���s"v�Tܚ�2"�uδ�<�|���!�]����<�qpQ��0�a�t�)�\q�[����,1���<K�Y��m��r#'IDm�����F7C&b��S���d��΁H>�	o�,=��}��5���Ux[x��V��l���/k�-ơ.;��gw�r6w"����k���a�0���F����;�&PӐUn���N\�(K�{���w��`v�����_�ס�]�H���6������$=lؐr� ��^�����uK�6�έ�7m����vU���T���!N����ƙ�Y�#ˡZ�����m.�UER�����6f0��Sв�@���2
���Ն�cބ�ۉ��-�zI�RZrge�xTb��X��o��{�����u���xaԜ#b���а3�,)h�+˄u֦�#i��z�Uǲ!�&�������ϖ;`5���T�r���0��r9��}��������G����Sa!
1�+�b�� �}�"�6U��(ٔ���#���\#�6+.]EӔ��26Ҟ��?ȉi=� �|���Fb�����E�-,(�k^��z��v1��=�, �K#� Gw�r[���H���{���|��v�ʹ��/B�tH��C�M�af��V ��ߺ��c)����2T�HM�&�A�{��G8���/;�/�����Fa��Y��W�O�<���ӱ�'M��`�����'�k�C�K�}�Os�S�����{��������+�Ku�H";��wD*� �۽Ԋ�\�$�WN��R��k����ShQ/��(�ٚp��$m����%vO�#�ji�c�����|h��3�����p�D��.�-��5#%,К�,C�8��߽���#�t�A棠��������E��w</Em���#��<F�! ��/�&p�lR+�e�Z�Hwz�������ޯ��������hqV�w�����f'3�C:K|�!&LN�u�����T����m8Ȩ$
�	3���b	z� �|���-�s��qp��s�3�XY�C����Wו��^��b̛����م��.�pg�c�m�%�!Y�{9�D�>��R!z�ɲhI3�͏��`FS;"�/f��ďI�F����N��֩8��bCRM�R�F�.�u��|�Lv*YR�{�*��۴>��d��a�3?��52���+@.��������l&!�0�}�0���ǻ�@Kˣ����H`s��~��:bi@�N;{~��-��,;�g�+�.vX��,ϰ������N�A��:�r�$t�?S'�z�1LUa������,���%�v:��֜V���[�>Hc�+r]U�g0Tn{760a;��Wݒ�+������aҙ��Y�L��JD����e��1-���Gq�Q��9�C�/?O�d��l�Ў���?�/K��Ԭ4~M���rJ� X�6H�V�Z)ο���y>R(�h���jڕq@&Jgp�Ç&����ڔr��i�I3� ���A.#K�l�����������i���/c�s�Ӊg�D��/�Dq�nx��tk~=!���a52�>W��k��8A����$���I��]��c��~���|j�",����P.�����J��9�px �T{���1%�԰j��pe	�.�$� �������j�@�P+�8L�%�)0�� ��O���X��t�n�F�CT��4�O�园.�H9��VBć�}����	Kw!_ l
3��ژ�n/y}�Fǎ�k>~��"�S���*��Ck�#"�Ic�����N*�����G�]��^xԨ�|lZ.��	��F�7�������LE(�����0��O� i�S/��y�5
��|ap�|�&�g����Ʋ�n���O}�sy��5�Z\���Xx
�ڀ�:IO�=g��]�Ns��]��ya���xй��/9���iq���6��K��\F��<���g{��@�f0u��e�@`��q?"l�=�lR��W���>#��n�f<ۙ�̰˳���7o�|��c��g��Tb�G���E�Q�����!�T��Q��	��
��u�IKuzt<��9"�V���փx=�J�����s����`74b�!�q�l�No֥\���9��P�0_��<��6��KB��ѐ��g��F��.���9{),�@��kZ�pJ�|Y��:ϕ�ܐ�����������U�a�`^Ce�k�Rl�(�F�X[3`�a��r���^����J���	 ��2v�vq1���f�|{8�������j�A����5��
�j�g�TR�XVL�\ʟ�8�i^�9�g5�Th���g(���� ����k=C���L��h��91*�B�l��<����w��W _�<#�p��꼚��:T2\���A}��t[�����~h�u�xD��6�r�x"5�9A.����Hvʫ9�d�zlO�dO��I�f�]}3�\�"�*�I//K�&�FsM����<��Ѭ.k�-du'(B�Z��G4pC��aQ�E����%3�v}�G��N@�Bo��/�Pw͒A�"��}��X��F_��x����%�ҟ���l���,S��uD�+���i����+�:��&x�>�]��D�
@5h�����U��~!�g�
�q�+u3%����଼��qU�o�9�����Y�?��Uy��!=VOm@e�|W����B ��<d�$9��X�h�$���,x� �49�ە�ͫ.�g���PKЃz�݈�A�+%��7�+Ҳq Ϝ��j���������2(\����E�KM�[�>EF���nعXs}�|6��"�斐f�Z&F�	�d��$VՓq^SV���28��Y��td+��A�:!қ~m�����}�E'�z��R�4v���f�ڙ�����C�Pe�|~5���C�S@��hbo�iU��퐕��!�r��4N��2d%�<�)!nfR��YB;��|,0��Ss)<�V�;��Nߴ�vlW��Kv́�}V����|��5���f��8�29����C�j�jr���<��A�0��	�=$��J�S��v!�Q!Ԙ�U0T<�'F��d&��Ry#
�����CC�q�|�q������ɷ�}S�'���{v�/ٚ��%U�ڢF���^��7Ϫ�q_P �
�.T=��qE7���z�R�'0י���Ԗkg�p`�^=��[���:��P?�v�Cl���4��8��i땠a]�Z���X������3�����BO���X#�篥��ߥ�'~A� �9� BZ��1=[��t�Y�W����mn�%�Җ���	^��<f<8���Ap㙘 �����H ��
�h���QHe��WK�k�-"$��)��+�ߌ�9P0K�8�����ZI�+����]ԂB��K��2ԌCGC�ﰩ�4��y�[S����gv���&޴n��e��n0��scC8k�#L���V�Ұ��@Z�R  c��Ο� ���� ��܈�J�l���$�Kc��p\�Lк���-:r�ׁh�wv8�+����k9��& �q1�->yB�~�+d���2�9Ⱥ���"U��F^�z��g��=�Xq��G��2O�m�~��E��Fb�u2�O�^~�q�n#0�}�AL.����_��ua&B����@WpH�}n��9�):NЅy��	����5:��FHϧ���$���"�3lL�������e�d���l�?�$+0m�} ������'�T����T������B�l,(=3=�l&�G_׌���{��6��_8!��@�����(J2Aw�x��K���w�����${�x��9]��c�nQ��7`	���J�D��4����C<%��g]�����7��2^�Q�?-M��R�5�*��jMW�٣�*�u[�>��,��x���N[�����b=�\5iS�W���,�< ����M�k�Q��Z��K�HU�\Hc#1�0:���?%���5�7��x�I�)c�{攥�6�'��yg�5a`������^�Sj4��Ƚ�l�%L��p�?�,�� ���KE�4��e�����"U���[D��j\G��6&�?��b����B�h:��Zl�$�����#��0 Y�����/[ZA�½?=?� �*�2^5^���K���;���������qGg^����`�p�Ļ51�ʢ&���m����}bfTO3S�E3�Gi����z�k�o=��D� ����.�ux*ǐ���{��M�H��`�Q
�@�����e��+�����hTf�o��Pa�zUԓC#��@�����=�{򾬸emd��S������;�u{���5�E�)����Ө8���9[iIĬ�s-�O�S����`�Mm?̰w�����a�.�E�38��s.h�R���A�|�˒}�U{��R�Ɔ`X�\ht��������*_�m��;w>�B�OW��Z��<�<Yz��7�P4��Rm[����|�d��Vj����B���}b��vfs�e�D\�0^�*e�q��-*#�m��o*��JK�Ү���A�����Ira�W0DS%��t���g"]���D7�OU����x+?�^,n;|֤��y�j�Qiwf�~/l2�ÞÙK�.] �>�!l��^�2�8&�I\�*��x�19��Ƞ�"�T�ڟ�-X!�!/�&�{~@�i�hG?�q�ӿ!A�'�����| �@�~�����¢W!���R��1ޙG*Q��?~���7T3ȯ��Xy��۰��E���Q��zA�%Ҫv�mX�_h�,�bF�����d�JО�E�^��ͥͻ�/{Ӛʢ���(�-��X�g�m<�`+C�V�`>+�oj�N�_� �,��H�Qx6��:�̦�m�����������rdV�Qu5F�&K��gGÕ"�����uivNV�n�t�4�U��<�E\�u�i�Pځ�N}�oxE2az�-P&fk"~lj���5� ��5l@���(ү��ވ�4��Z3���y��ڽ�Y�Ɋb��vޕ������hϖ��Z����<3{��9ޥ31���]�/��ٍnAWaQ�J%�@~���XJ����b�%�:���PX���/[��2�S�F�T�|D�ٗ4��I��0r`�\%z��ĴZxT��rus�|ߒ�ɢ��'p�Um14l�oȫ3�%��,ط�M��B�OЂV���H�x=�2B��I��܀�8C$:�Pk��`��:��'�s���b��.�	�-�#�� +�y�:���O|c{g�͙w4a�n�T?�?������_�u5m�i�e�fQ�<�[!���Ǫ�XQ�k�2����"~x�P�g����|x�Dh�{0f03��S� G5p>v"�Hjge"��YV�d���(��M��=���t)�CܐU�k�7�oD¬��N�{N[9�^�g��n��A�P�K��-c�Q��@���ٯ)me4nԾL'.�߲��)�a��T�)�/�w�,�>�V���,����{:v2�q��:���'p�oE5���P��>q����7Q��-�.�y��}~��Zj8���<a6P
�'ag�,��4"�J>b�>Kӊ�����jTï�hƟƊac�*�����l� EVJ����j�P�����n#�@�qT���A��I܊�ǒ��*LS����_�LU��5��7|{<��`C{K �ߎ�Ea_��Ok9�e�e!�kA�|�<_���h�ܚn��8�ts�\M��[���+�=�	M��X9���ZCT�f�H~V���T'�|3�"Q^�b�9(�Ch=�w�nhH��������S2��g)���%f�!�m𥌤Q��R����QP��A�OHQ��2��jv�*�,t�v�׼�4�S�d��X�b������:�Zż������^GLI�e����Qz�6ę�x%'1��nъ�ϯA��N�a�BI��B0�{܅ 8��8���l�V�o��C1|/���$3ꎀ�����@�{d��������9^l�Q�q�j3������H�V�R
 3�������ꮐ|�j���O6����������ihTp�$�i�4��ƽ�T���eo~��wr�?����8q*@v��țkr��|$gd��ow�X��☠W��\���a�(���n'k~��pP���D��.aU��w��dO�e����b>��S�sQY���w�+����t��ZA�;��{�0��`���Wq�I
�q-�_�+5�/�P�����{z��O;�����~-3�O6gJ�`�i�]�w�0*���DLuٞ�y�=`�}_O�(���&���y Є�]U3,�m;�@F��Z{߮ ]�w1��� W�H:l:��?u&��x����)���{��Kd��q��Ua��Kl�?t�9iMG�J*�1��1I U3�_ �>�FN�!f����oxRF�/A}<���o&� lb��X�0T0�f��8��sRB�ej�2Y �S�R�+<��&	XE`�,��V��������;."�z����2���It)d���ɨ5S�]�����u ��ÍB���ʼS��ޕw�[��T^O�oL0Zb[J�"�َ���лM������V��s�'v��{PpKR|�XV
��$�8�Mn���l��$C�J��Ŷ������K9����ƨ��#y��?%�Zt����.���w2��奄)��$����-����Q'�]cM��!�e%����nW�b��Nzh��M��ߗ�z���5��u@�����;�;K�+#C����	�tE6bI �����yٯ� �>S;�-z5�����T7��� ��`�2r����!`���
�E�f{K�M#�.�Tǔ�C��]I��Ad��	2��A�C8.�'щq��|�6�Cfl��uT'���aH���;�5����4l!e�`D���	���ebw��=�0��<کE�;\Q$Y2/�'A8��~������8��%yq^�`�tjuR�i��U�p�J��6K��Z"썃����e���x��(s��4�z.n�]�~_���gp��&=���`oq��a1�PaKo�����(/��
�sY�)���+�����x��KN��������M_e�g�8�C�W�;�'��]Y���P��%s��%,1?0w̞`_pJm����T���K��]�"�@���E)��#�S��ڔc��Qmq�nQ|���ia��ݛ��>,�4~�pV�:L�*��#�=iC}�`�Wў'AZ�1�Cr����Yfx�)�o���ko8���F݈�=�H�B=z�_$��%yW_��_�B�f�XM���9��o[��8.F������jΛfޗ8A\�*�"{���{��lY�]\���A���q�@+أ�s�yFwA)�#c���&�w� �/�W�3�NR>��,Rb;��
�h��p���g3�b��\����e���LZ��(����]�����(�ޜQ˰��PU6e�[ͫGsc��+�'5�%o����b�H���J�:敿RK����j�A�m/zP ��La<<
�J�&�R�x枣3�s��[�����S5�S�G\�y�f�>]hn(�@9��5�h�Sk��)��p}�\��X�k3�?�r��vto�/�����@�`�C�y��D��J�p0�(�j'���N�;�BoD���tZ�.\|�y��������:�Z`��S���H�p�:�ΨT?�
8�z�-T6��Z��n��ݳ��Ѿۉ��?���N=	=��xٱ�a�L���?����ĺ�h�[�NL4�捠�glK1���<�����&n)�	d0-V��T�[n[]Ǥ�juۿ������*~A��jc�Bg���Aӳ	mM�4~K��V'�$�'�����ર��U�()]��~t�@�u�}}���3��?�;3`5�[L�H��%��ᅉ�⮞�?_n���ߒ��F]X�(�F��|($�ϼ����'ҞsB)����%,�yw��Mfn
��"F5��A�bh�;�t+�69$����o��2����SC7-LD��=b���(�?��*��lFAՓ*B7BW�_yl*��?ͤ�iݸًcv����g����6������/���^���į���33�<N0�r��G,�ȡ=eT�e�#��O� ץ�����'�?����]�q�F��^��+j>7���w�� �w`W������kW�#TP`��&�Xd�\YF!��ޥ����'��K��RZ��o=U����XK�[gZ!T���ob6�C��)�jO��*O�����\�q<�ԚT�Q��a��(�V�#YD �x.��/3�\)��݆4KJhi�����h�ari��~`�5��Jb�2�#����)A��g|C�ٮ é0Xť�ol��A0ʎM�$����e��6�o����`[vg��/� R����v�.��I��� �3_�_�:���ٝ˔�r�쥡����!k������>�d�{��o���y�ßI�=N��B�z����\�h���|��o�&Y^r����ոބ�N�@�t %���z�:��W�6i�Tf�K��?Ӈz�2���c�f��L��J,-u矾���4�?h$���D �.�1��<ck�>1�P��B���IDSj!<v�&�`�`�V���3�[Ƅ)IpV�$(����#,�ڴh����۴�Э�AD��L�։~�`˳;�W���'m���n�S�Yz�,��˂���Z�
��98|�l��h�ݻm3�|}������_���(Ձ�嘊\�?�Ҋ��C��p~��A�I�^EH�5)�.���$4���,�D����)pz�e���O/�� 闑=a�Bm�nA�4�����v �.g2L�(/�1�>�Aj�	��zŬ(C� �	�5�C����2h�UD�@�l�=�����^�ӈ�W�=��{1�	�*Qt�M
��*��b��&�#aܨ1��M��֯k	�f�m�!!2��c�p�[�c��|>:���poFm�o2	�~��¬�Մ&���R�HCє2��D�$��d�}���"qɗ����tUC^�)�N�@J����C�k�H.V$0A=֘ፙ�@��~�U�qgw���v+4 ��>^+_���5�.�84?�����/�p�|`��2/+�*�Vr,�2���hR�u�� ��Q2��o�Rs��M,Wjrl=﹆C��'_�����uЛ�<o���uv�?=)D�q��I�\GMF�h���y�vEG�R�v��H�=����4�G2C��B���b�����"
|$t��LE �i)�vZ����?r�"�o�ƣ{��m�8_5� \���{n\����^SGve5l��Q�E�l��F�;���j�6�yAܚ���G�>5$w�=Wl�8#-�Ӗ(�� � (�$������ͼ�$w����H�/Z�<��]L�H�ei�cfܶ�)ڙ7u��70,`���/�����:^G,'\;�[R��T���̺��|���ޫ�K�V�yV����.��k��W��{gߡ>��{v̫1�ڣ�ӆ�ڞ��n�F�����}�0�ؖYG��w;ϱ���{�|܍=՟�t­�	�K~FKˊ��(GfM�H��I�V xFz���q)���N{�9�{^�m�?�M"lSX�j�Đ{����nC�i�k�l!Qʍ
�Ah��`���+k�<�
��9����Zgo9L?@��$B���nC8�1��6}�t)��;��.Q�G?��hE����JzM�Xz¸ߝw�vwB'���Z\`t����1�ĸ&�ؾ�c����Xf��ZMu ˤWo"�
���
lh�� T�]Eh"xd�f��0���l�3�T���mMh��?�,����*�e�K⶘I� �g�&4��\;�?��3�*��c����ur��jP���/$�0��r+���i�9��£,ﰝA���L"O}�P��G���A2�6��gU)�(����2��ڊ�����S�C�*,�G�����/����yM��I�M�E�q��0�m�`��G0t��/�\�vv/��w�N���9H��W驻M��\NP��k�s\�]����#�تŵ/��@D���Q�3ZB�Z2�:|#d.�C�n���Vi��.�21���9�
��8����������x��QB�)0/V�*t8}M�8�Y%�tVc��+m����MM+�#��%ӎʉ��O������CW�g@Xt���?em�qv*#M�������WU`��\]*�ҽ�	z٨�m�ӏ?Cx�w�!�,G���y���Lp�{F��	��7�R�7������ o?��{Mh�:�������:k��Z���BXLX�R.=�~:��g(�H�V����M��\��3��y"��]��݃|�z��$C���5:�����U:�l�ڑ�G�5�R?��0�"�4Mg�Ԑs�-���}��(+�L��aC��o&���n5˟��$��r��5�D��t���vk����.)��L+=�H��6�DY��(O�"����!��g��^�c}w:�k` �Irzb/�Y�d������
��s��ݸ'J,�B���	%~���`�ae��/�ޔ:Y��eM�\2�l͔E`��Ї��<NP1�IwC ��TO�u�|+���k�ͽ��@kwQ�={9�gZ��,��|zfjU��A�&ϖ��\ų��uUʘ �۾[�'���%<0��\2�%a�̱:}4,E��O��م�S�?DQoqf�Dxq �/-�cK�J�(��*����D���Vt�`���`&N�Kݚ�����,����*#�+����t��7'��R�]dl�@n�#;g�����8x:��_@W���e��p�P��m8[6�h�ߢ�Z�Az}�[/�`'���&��y��}��Y���}Rj��g1����rz��%q��� /&_���,�Q�;,O��.:ݎ`0o���(%�V�?S#.�BF�����J��_x3Z�`�Tn��d	o�����d�4}>c��0���Ge�)[RN�3j�g��+�+�~�U�U��R_�
�S����X`5GGt����5�bz���{�.Q'�>��<�D����Is���x|�́�P��4�%%�p�|�U>�0���v�95�b'�/�/�	�rmO���Q���wz��f��^�0�;u�׿Y����	���56��y��k����A���
$3�����l�CX�3{�4�NP�C1�]L�8C����y��:�ݴ�6�P��.���s�CJ������#'#� Qg�wOY78W!��.�Od৵R�d��ܙ�1���:V�ˏ�L�Hġ\pS��V3T3�!�<�/�f���?1ע\�$�Y=���~TP��e���jx��,�9V��zzL�P!P(�aГ3f��7v���ha%-�8����B��	�;h.�`�k�G`^���2�vB�n��.�Ang�����8��"q�M��L�xF�����?y��%`&�n�W*�^�5g�����8s�Jl����L�L��ַ|�_��q�w���1j�p���2���<��[��+�S�?A�����5��9����)*�Ҡ Z!k��Y�=|p�,�~�K3����t΀�ƫն���'C��� �!/�k�_ 6	�Vu.�t�X]����Z�S�;|D>T��a#�����=��o���,T7��Q��=��ԶʼD"�B�����-�B�24��f%P�E��4-�*�Ί�����5��JI�]���0���%pC�Y����q�J9�0�O(5]��p�_ [�s;%�c����+�A@����؉�g{�ң��ҭ�������2$A$S�,�=�D����=eN�rP��-S�n����=���$I����O8;�V�2�
;�q[K۸�i���u-����jћ�jJ'�Kx[�N����οOaX�FdhۇI(8C��o3����?�D\�(c>�ͬ��!�ג��L�h�~�8��#!�(_,,��Ս�0������qޟJX���I�[��tIq�(����6)(W��F;�pY�T=���9z��֮7�ݒQ!�T���:��%����,�z�����[pi�������	�����.����敯��*Z;�&A?�q�(N��� N������Ƴ��b�(z��6�d�ɕZ�H�C-���|~�L�$�wV�#��'��4�	��\c�$��\~���t"K?OKt�0!�9@YL�Ö֟��?moX/��υ�j4�;��@������~q�5�LJ��L��%��rGz^;:��) �BN>g�O^�R�f�]|<qu�����`�� �
��u��_p�~�>�����2�s.��cV%@�P]�5Ոv�L�|��� 
g~P��<)5D��g &v��=��\���j��KaY}7�w?�����Q���ʢ����%W� ؒ6����<l0��� J��b�s�>��=�VP,
����oz�P�K�����*���y�RjDU�$�1��=׆O�ra��4xb�ZŜ���)��+��W��o�в�4�[�:���~K����K)�4I|jݠ�ֈJl([�� �$͠k�o�L[���8h�"��d_Z�8hu�	__��[l������%�I�[b�nv�k�xu�����j��v/������JH���L�E�\��T�OH��SQ�������͔y@*N��!Z�m��@vD�'=��ʺ�������'޶����&�e��аl�g�^�[9~�v���K��;^Rt'l�m����i��  �e�c51;��ͻ\��i���+���Ѱ~dډG'",`��b�X���(|���Y�c�#v�h����ݦ�4A\�9=YѤ��?J|M
��xs�7~��e��Â�K/�c;�۲�y��~2��=�Jn꘧_}=w�;h��Pp���S˫o="�K��C���8�����W�0 ռ���Vxvgt^RjPEyVdtD?S��K}�����}�@��H� ��r����X�iv���ʡ)U_+Y)הHߵ�V��v�����%���٧C���|�kߕ��=T�H,˛c0�.w	4I-�q˶���Y�f@xF1V�.φ�D�e��Th� z:WJ��������������j��O^D�2�ُ���[���2��=�X�0�����q�e��� l�0��ʀ:���~ArmX�b�����Sp�9���gL&�l^ױ���n�I�FP��hX����a�e� �I����͔���ջ�	�aW2����twہ��@M&�J�� ���b/�GM_e;���e'_���C�����o)��/hؕk�/��������[p�7q� /�(ć-���vh�#=��2���$�|1��f�V�?�k.�� ��x�G��)����a�6{Jk��36~�|���]2m"��~��+�}b��Sc~^�5�:�E4V\m`)���s�ɰ��#`f27|�B�Y�}_�7��C�:��y�<�����3�7����!/�ݪ�"�ʭ���Y=�4`�L��ި����X������k(������o�YމS����eus*1�ժ9dv��<'(�։0�)�9"zQg�\�.���/��\�Z����!(=QD�v�S�Sǌ��x�Bq�?Y2��1��$�I�s�7�=-n��}r��|e6$Ty�\4�y�T�VW�K�&D��@�W��b9$�I*�	qvp�:���Y�v����i��o��Zv��ϧ��v�h�z'i+�s~
��������Ë��N9c[V�f��@��2���*׶g�]�	8��-�n[�6$~IC9vu�I&���g6���. θ�>R95�tC^�X����GQ�Δ�H6�`��C71G_� �U�<�����hv d ��̟L%��v ��Ge� �RE�cvaJ������!���hY����hb��rR[�zPo)��Y����,+\lWsda�5�?��f�=p�6Wn�F���)�|,� ,�:M����/1�%���0��Lp��riZ��HG�Z�S(�!|	n����I#��TR�]8�CckĊ}N}:"	�oft�mӻ�
'�~J�]x�*dU�·�2u���[ưe�#8|��az&7��K�T��꒠W�쐞7��9k�z�[y��9�-`/���c�펟���9y:�D�Gʈ�]yԇ��oƃ�+w�hB���3��u ^$]T��PGL���� 6�ݍ����sq$9�t�*ǎZ4?"�����'���_�LM%g�ϊ3�
l�{9��u߰DhΦ4�_i}P�䆂@Q�������z*�o�;���/뿝��i�	O�3�GRL��k���F�(�i��FKV�����K�����a�
��ց*�Q]E��B�{����B�߯�%Ծ1�`��ҍe*�g5'[��Q�l�*�L��p%�@=ז��;�����z�'��(f�� ��IE��^��
9�.�b碤<��m��\��g�"JQ�����܌l,)X�/�C�>[p &�vz��vA�_��S���9@ǨX�2�����gp-M��L��w�L��K�ߖR|�� ��]j-��͖�}B�w���64ֆy.�k(I+��&NAB��Z��u�����YMāz�����e�*�j�v�p""��L>�E׸]e
r,>��Vud7xp��˘%�N]qb2Y,w���e/���Ǩf�U�x�\7'8=�7����?�$���	�A���~�	C�u��l�w0�d�U�y����@)A�oĆxA�m��|�DPT]�� �ld�um��.���`虴0a$�B]�U�ۂ'�:�^��|�&J,������)Q"���t�R��H�*�����+@�휋@��c�Ja6kɫ"�\oY���h1�PLt�z}Q����	���6̓9ז�g�H��aٖ���)�f�&�D �V�_]�M�'I �҅��j��#K�8�iFﴪO Q�m- ��h���{������$��,�A�ӥ-�:a������_N}8ʜ
[M9)�T0	�B���.�q|�=t�`	�b����z�%��~?�#�8,�o��S�Y�18���=	*�2av�|�e��ǿ�m�pV�
������b~[�m��b�9:�@��ab�o:�^�i�Wݧ�]���5��o���K�q��*ؔx~u�����iL	��|MA��P_Ǿ�BX��p�}]MM>WE��q�5!�Ж[ "I�sg��C��y;�HP������a硺�#_3�B�U���h[c�v���@�b�$���Ƭ���F��ڊ;E�������u�k\̐yU �a�!z�������Ԅ���;s\9;3p"�:�
f�\���S��cz��A�i���CD0r�(���N�F�FJ,R��n���֨�3E�m��*��c����|��dk��Oٸ)�(���eΔJ-��Ɨ��tx8��#����&N*��F�J�uǷ1����my�ڎ���a��R��J���FA����D����kn�c�����+�fw�$�zZn,���&���ܯV��E�������ڣ���@y���'�u�@X�!�Q]�`���w�_�9����E�]N�g��D~��!�L�q�V��PR ~�~��z��9+�l�|L�-1;Q�g*�s��t1u���� ���ʷ�LuF�A�l�+���r"���2>E��9�Ko �����Mث���.��{����(ǎ��1<<҅=�옥�?Y�&F����8����M��G@J����-��᧯M�30����$���&�TéD?s����]�_�	+l�_Y]g�L���;g�������Tl=W,T�'��0v�35� ��E:��cqBd��d���P ���7��5<�Ͼ�%Kv�uT�3����1w_��M��o��w��l���=>{^������{�H".Y<���b�hϸk�D���oJM��ih�"`�D���I��,|6�o�$Y�K�f>��Ls,��撝{�P�M�s��)1���r�k�S����O��`<���8?73w:��7�ӝGP�t�W�S�S�Q2fx+���$:���l�>t�N�^�tʨO��]����s%-�]�̺P�R��ix �Xo <�z�s+#VTG��VF�P���]|��ĎX��x0,��Ǐ��w�ႋX����U���#�
07h��8��V'�h��]�2�2y�:%}Ɍ��xk�Rc��m9�6ơ��N�+�>�Ek:W�щ�v)>�j�'d�xE5Ԡ �ȌC�1f$�Y�[UY�0Bɐ�����4b�z�a��k�+f�^kF�O+AG�Ζ�;a��«()�2��m6�HZ��!���i�{�Ӡ�;}'�H32�R��&F])jă��2v�A`&3i�k/;6�����r���*�Ƈ
��8j�9���j�4L��n����,߳�Mߛ�Rv =�M�~	�zt��`R�4�=C���1�e�t����҄IH�w�者`�"�$�Y���.���Kы�������k�9�W���?nG����j��Mw�3\n���/	g��.,��s�C�*5W��$0��ɦǙm$������U�,��"���N0��x���:%Rm�C�Y����r/�"'*�7�pK��E`�ܜ}�4t*8�^���H7�+4t�j4��ywW��T��_⏷Y�Wٹ�@�5�Rzt��V&,��hBUR������;��+�pv�a���N���ĔYMs�	�7ލ&򉹡�K��%�!�������e��}l�6��*�*��ũy������4�>g=�X���.�ӍK�ju�*{�8γr�Z�5�gD�� �˜7�45x��D�#5G���T��8a4'YO0ԾOK�4�CR}�h�A���B8(w���� �-j�F�M4]׫Y4��E����j����� 요�F�;[H��1i㛻���1��������)��Dܐ�s��(���[8g�tDgn@�u���X��ؚpx�i�������iώB�>�걸T�3��Y��x�U�]��f7K&�	?1�z���3��V̍a^��<s����n���0Gy��	=9�φ�kŶ���'!n��N�������mN(D��9��}W��\. ��Ê�����jمUճ��R΀��t��=�$՘��I댜o ��xP]ZЗ��N�D�g��3�ј�Xa��U�!-w���}Z� F�>������j���m��%jL��Ey��v�C9�W�Xd�!�4 �v�#C}���uO>�QT3���-�
&�fe��?%"y���q�5BeWV;�gx����J�iU{�7J�(��g�70_%�6| 0y�%� H&k�j�`r�/l�u��Mi��	!3|��&H������[h,����<��Y���̥-3���Ӂ��_�#ySUY܁�so��R��U�b92�
�yE^I�q�p"tԏ�jR7O�ȥ'�����
�N�4���k��	�d��o�~_8"	��f(��U��^�k�	�~ ��;���\S@��m��r8���0�\/E5|�����Z�
��Ȭ�'�:z<�'a[ Cf�
��46���>�M&if�.�L���>@2D�׭^��9�̗���U�z.�@��vLI/k:]�+K�M�̻ESޗ����P�gH2�����ĎN�-���/�i�R�I�oZ�G�|����Mh�T4��
��Z�c�mj܀�<L1�eH��'I5-R�TՄ����b�1F+!�Ъhd��5���We��1~"������.��혅��o�܊N,�����Uvھ����Eg���b�ydf��݀!Y1Y�v?�?b��N���x���H�"?�z��E6H�|H�jɻ�AL��@�f;��\_�;���c����^	���v����I����(4x�P����N�"M?4����L����~M%\�1���!8��G�4�f��^��!�~��s�,6,zh��_W0I���9��c.ZHȄ���=���Ĭ��E�rQ�bw�T�6�ġT�1�N�4l��V��Ou��԰�U 1e�8�`����wL�p����h�s�$T�����cC��Zp�p��9���陒N:&� �x��z�L�V~�檫�>2�E�����,C7�4�U��$��"@��x��7Ev����=��̻��fIB�z�V�Pi��1�1���:&I�j���@��p�`q���Y�v:}�@��n��RK���=�=cA�����{6)�������i��@��ߙ�+Ǟ�W����]� � j`,G�#u�|#��f91)��)(��Г:��q,�0/p���4��S;��(����ż莾 ;�w��7@��l����o�	�x�f#:��ۆ%����^�L�`?s��.�w!��0�_��\5i��5���
\���vp� [�GgCRe�����؄�A��Y�L�%.��ܢ�����,b�7���qߞ��a�:�����������f��:q� �"���D�$���qHHE��K�|0�Zl���� �N��A��ve�/-6˗p����F�]��?�gX� ��zfj3
�@����.�sɯ9p �e�B�Hل�w��u���ڙfё��C�m�-���{��Z\�|�e��Wm6ة8u �07-R���3���1S�q�O��q��c��יɂB�X�53�-���HA��2�x�?�sb #_L����;��͕�ӫ
�m"LO:?@}-�����W��$�#y����*�5�`�EB����>wf�#�lx#��@�٣�ƶ�'�Q�k�^r�\3��"2W�S�_pB�w8bՀP�*)rB.*~lp16�wS��o6�pS�S&3!�χ��e[�$�n_ٲ������@��4�"R�0�@�Ȧ���m/eVɷ����`:�,��s�r�ͫ_i�$bj�QF.��������奸���\~�3��t"I5�K�s� i�����V��1��kG/Ң�PCT�GAl�ճ\1䙥M-�Sv<�:yq�W�{-w����g4��]�?ܘe,��mLA����Dl��ḵY��݁��8�h��4#��\<x�'<~U����CƪVl�r�Wt=���M��6	;�Yc�ւ��O����-��._���@�������G���x�|}s���>�-����`��w��Cf�/�
�T틨����3�b��Y�P`~�+N-��� �h�V�k��~��0 ���������^���z�Wx1�Z���8N}Ր��'��b{���LgH�����$)���f+��B�}���Olf4��b-����8�q��a5����+�[�a�g��6W���!�K9�������mHK!8CrM���ԝ_H�+j�t�[�MD��+�ܯt�t���c�`��`� ���zzc��v��Z�;���tV��Jꯀ%GSTy��Vv�[q���j���i��w��_wEl�z'���ӆ������<�QR�4W$�����!޾0�7��r��l�R��S���EP�<ځG�Q>�����[zDx�w8�S�������ga��+���[ub�� ،��\g�ۺI� >�����N�BI������I���^�̇�I6E;G��˰��� ���2p��e�WD_�Ȫ���3�5Z�+�F�dJ�Ρt���6�4���5<z��j3��-��H��.���WA�[@Ӷ�C������#m�_L+u�Zk{5�^ڛ��FAIww���7���'<�pP�֖��h�\�����MfC�G\�u2RG�2�Z֘��,�>o��q�x�G��4�HB� h�� f�_ǔ��m���(k���|����H<�zr^���=���c��&�S�)Z�V*Y�o�c4{���vnFg�4�8�������^%�O���`D���iY�i`��~ը�7Shi��}� �O���kR�E���gk����HP�/��a�~`L���:�I �1�E:�ȩy��
�B��5[�q*��3�9<�wD=DfR�`�S���&����M��=�<�!��H׫j}"����a�s��+��Ɉwj9��H��B��3�#�X�~(�uD;�".n����z�ǃ�20������73���������B�15�2�������D��!C)�}%{l%��4�b�9 Q3(�S!�<YW�j�����U�ƎG�`���P^��t� �S�ׇL�BB��0	W��:�6��n_Q�h#Z��,+���Q�}żw}��Q��ڎ�:��N�ϖ򪊵f�`3�>5\Va?�
F��m,ç������
�65SUV�K�+���T�Ed�+<$�����
F%
�ɰ����� e����Ij���G�aBHԔ��T���d�3K��E�+4O23;�(B~���ۡԋ��Ǡ��j�3�o�Q��!QMVOԾbX�� �[Eg�Sd�'x�O�p74q�9W�2�<��M	ѧ`�F�f����8���' �k��cS�Zje�1�ںa5�#��Ww����*�<T�M
�Cj���?x�>�`3F�~��5
����6�
�l����c��^��Ȕ���)c�t�;�f��nz������ԧ���ݡP�X�B�æ-*Cޅ-�����.��yH�:7�D�K���叏��O��Ig���p���*�ؤ��9�s?���M�(�Qh�f`҃.���\4�z�V��ȏ�
Ѓ�a�J�>��!E��{OO��_���Q��A"��P=������I�����j�È�`X7Pp���OJ'j��!x��� � d�p�MG	�J������ĕ�E��$�,�๣'�>s� ŏs���5�T�-��R޻̵��q��ѽxy�:N��.eT�?�D��D��AB�3���ͼ�����wSŐ�6�*�E�6^��/N9 ����w3vٜ��|���w��)�x�_�R_u��sP�@�MV��3$��-�+��9��eyG�v����!�O�N�#-���2~g�,G�������N�~׏v�[��kV�z�,QrtXG�"����;I�&h��-�@<��/RS�лg��N*,E��Y`M@�=rFc�l����*L��8�H�!�Q���*�'&O�%+�EI�v��}���x��bU����m�A�
1�n�xp�e��w������z�*��S$�W�OȭoTF����Iƈ�E�����(�w�}��9���jЍ��MS���P�[-��֓f�����H�Q�h��ع��G�I2���:�+�f�n����sø�"�d�����������N��o�֛A�@9��B&4��;	󿪛l�������,˞��N���5��d̖]2$ ��Z7��3�����[ް��!�O�x+a�Os(�y8Ս�e�~�%��(���[�2�\��@��I����K�{�H9�{-Ytx���XI�6\��`�(��T�Ņf�.�]Pk��rB��~GY���R����&��Dc؏R�rՄ�	A�	�3��m'�G?��7�N��(�U��������)�齇D��U�X~��u΁��N'�����.��� j�)Z��ք��������z�����&P�� �Y|�)V<��%�o���C�An�|*]�/�r6Sw�!����<���;�$���Rd�!{�t��a�����#���t�����ߍc��vͷ�o�Q{� O�23�>#�jx��cy)��,bfߠ�3�D�
�!
S��FkE�3���<�/d�<[����ӷ��&t�7�+����5�2�]��+�4DhrE�d������NJ-�Ox&0�h�(�ch��^9w{Rh��o�[��?�w���`�ǚݯ�/Kl�yV!��q��ed�g�
�*l@o~pL�ե��a����y�#(0�W3��<�D�#el&���zV{�S��~��]]�t7��[W4[v��z�_o,د���'-�(`!r�]4 �p����д��5�!M�����Ξ�9�|�ϰ.ko^�N@�Z^�;�|'Z��;פx�+7i@��"��*�@Aq���M���Z^�@���̯Ђ����Gk�yv�>C	3�siv���Y>�Y�M����0���3��A
�E�(m�xz�J 3�s������T��\�a�Y����o6u�S����o+��Fz��V�x�L� ᅒ����{�.���Wӷ�a�ޔ͝���8_��&�k�an���P��$[�@d��`NQ,H�i����|�;��(X�������]��7�n�P��{ٺ�_����)���Ʒ���k,��"M��k\B)�Z����*��Gȡ�Y6��)u���%�	�ކV#l��^s���Wy��8q{8�����'Q3ͯ&�mGĈ�Jp-b.*��;_�h)u7�~wD��vZ�}�sQ�fAl�-��7U?��x��^��e? '"Z7-��8��S����xb���cY�  �����?�Ta,�s��u��礧�I�k���_�<�Q�!5� p�7'0_ۘ��8x8XƚV���㴏���
��2�8Z�:X�"��ol�N4%����iw�i�[�����.�@8�`l��=��R�v�� "��D��m>��Ҕ��S�L�F�p�kҌ��a�Ϋ&�,�,�����r�Z�O|f`bT:�m�1]�c��g�=�z-έ\�B�9��+�bK��=�)	O���	\�Z1����ug��tB��I"0;�
3�0H�����6şn�b�fL_�)X}��Z5?��}
Y1y��A෉��J����PS�=�g�5*lU
�1�����Z�>��H{-*8Q����#����y� <ٜ�ߜk�b�E�UW��ee��6�U��55��2|�E-L&�`����4d!��ȝal��qa5X��S)���w�&�NZl8����Љڧ�u.3��M�O�&X�TZ6��~�������&�5@S�67��ĩ�9$V�cpt�ͱ������,k'dôXZ�C�3RHW&Yؽ	N:Lw�R��
�i���0�ri~#v�)cgJ�|DN�W#�; T�Pґ �z8�-�߸���P�ul��^	@�?�g��<Ŗ8̤A\�׾e�m��g9}(��,Gf���C>S�������83�ԭF6�S��.AM�8�"�6H�b������k��jc����+���Y#;H�\�2�y3a$�t���tN���h��%��C��~��	 ��^X=��Ry3{�*��z��U9�֘@Y7�у�¸��R������v��k��xA�#uӂ�#_��I�\�]�UG3�zj�u*@骬PCԭ�d@㙺�1���D~��'/M��G�KOm����F�ϰ��Gk�e`|�o։���Kښ[z�dT� T�1�vg'n������U��Xej�W�3�,j?���ZG0�Y� 7C;��]5�j�1P�td\� �㰂�D���ۢ�/%��Z$��(`�
���˂%��0�	�D�[�yC���n/�D��}�[�$ `����HR����"����DL���+عp��.6.wҞdVR3�*|�XV^ظ2<��T��0Cu��u�	w	�P�2sU��
}��*H��C�S����#�@�\~$����_T�7��8Ԡ��A=р2-m�s�ud��i>5��h��B�<Z�TE�	�~^�됟w�~��C* Ȩ@H��÷�&F�T\z�.�x��5���ϟQ*�|���ňk����ܱ�'�A�ͻ�_�s���tna�d�Jv�a�B�O��U���v�h=�Dֻ���{���� �-�E�|yR�9��ǃ��� ۾\~vvS��vZFö��s��{�^��H��t��@���wY�>,g�V�� ���Ϡ}3�j[����b��� �pjT��ih؇f��5Ԙ�!����A�ͩ@�&�Q�yg�Iu2�����ل[r��lH&%����t������o��"�L�q^3A� �3"�����!�,3������;�M�:��C1�m�U�f�1 !�h����w,Mn�0Z^+%-�t�e�|�¡�x�~e4��faۻ�ʖ���o�~8ow�SF�"?�c��G\m�`7�O���}���/�A��7#ec���B�&�u���HK`+�/t���U�94
��g�yM�?������S� ���@j�S��N�	Q�<8*8%_\��ѵ%� �v�gHݢ�c���9h��(�HH�JE^+M
Xh�7ހ�-��ɸ�AH����4Y
�)xA�}�0\x�:v��k����b@��GU�Y�gV�&�=M�pA%�TU�����#�C�ԁ^n�c�����͵������N�)���ῇ�Rq�;+d��
���ޫ�x�s�vxq�iT� I�0�/9�>�A�1�f能(���r�����< ��ϣ���v���%�� e�e�&�`l�G7��y��B�}���ʏ��/�C�L�fH{���dn�X[b�C�1�l�!zmb��u	�Ex�Y>3��pC�?�޼���o]�V��st.�8��\��;���FG��u�G��P�^^43Ty�1u.H�g!u��]�~�����e*>��{.��4�S�}���K�h	^�I��i/ao2���d�Bu���u�?�W3:��J�qN?'�ri_7�9J*��x�m0^-/���6���#�?�����3Fa�c���(�N�LŕW�f/B��o_�咣6�w�4g�Ȁ�A.\MX|e���9��)O/Jz����Nj���ns���
n7�+`aJ����/�o�&\Z�1����D�ۿ/A/1�,݊*�3P\��5ҹ���˙\������5Y��QU�z���j�$Z"F���w0���,FT�,O�_$������ݞ0
��12��:g�At	��wJU �C?�L]S������ ��$��2�A3����(�8\γ�PYl[���B�l�i������G$9í�u��t�zO����4�����%ׄu'sCO�g\Ivz/����U����ڃ����n�Kq�H�9d'�� �"�u�P5�9�,J+�I֕rɸ�NMR�nA�r��$!�����mvJ7zl��g�� 1�;��osȟ��(ċ̈.	�/z	k3���qH�n��%�X��h���[|�M���#Q4(/��س�N,����Wa5OZ(���w'���TV<�I��]����0�ɔo֒2I�~Z���L^�"��ɗp��F|ƁŤV��1u�SϪ����ؘ��D3��Ä�;~��"��Ӿ�Ϟ �R�P�j���+p�9yN�'�<�\�W��EB
�z�*Ҽ�V����f�vz�AE�U�Q��j�|?梌��csi}cxǑ����Ny�����I������	�`ː�a�ca�J՟��yb�<zZOQ�vm�n뇖{e���0�n�;vʨ�0��s�06��osYV��g�����IjYmS�	�����0'�q+�<wv`s���Ǖ�r��E���6��q>��%���B�#���C�u�
~QU�CqC��w�HL��b��NR\# 6l$����]װ(�`]G&/.��9&�54����`��p�7�7��|p�r������Yw���a6��tʱT�f}���Uz�x&�W;zx*f��KZ��tڠ�o"R�o����$����-T�edM,ސ����49�Q4��=��pn]��,��ϭ��������fA���:��&/u��%�
�,//-T�x�q 7i(�4��ȭ�����X))��g���jW3y$��4U�?�o�c�8����0d�bp��n@�h:���K��z�����3p��,��̿������U��-kC'b�>�[�<~��><䈕e-ܭ�n%?r�!w��-ߛ"��P�Gt����߅�2匟�����ȸ���8���N�l\�av�#�������qT��y�Ug6������K��,��rz�:su|.].d�'/s>h�G��/ Z��:�3MT���ϧ���z���S�+�mſ+H�^\��Z���V�=CF��)�︌Eq|㙽5ȓ��D�#FuoD��z�6 9�"��w&��c��}�r!4��)�"�gL4;�-��*؀c	�t�m>���[Ôr;N����eӫG'p���������'꟱��`�OI��ˁ��r%�$TQ՚�Z������^��|���t�]ZXyFc��uGx�r�h6�E4R�!���D��
yg��AdKB�^]�;y�/|�R�<�6�O������cw�i\b&{��h5�[`�iG�Oũ%�l,+=.C�Bcճ�{;�!�S��v��6�X��WK�!�~���-�W�;3O�O3���S/��N�Z>�X�v7�1V��2Q��$��Sal�v�].�6lZ"I�e�ņ�&v>Ͻ�M��M`��(Bo�ՂR��>x~�XAl+�k��P�O�3��*@+�3%%ʫؘ�1��^���@���k<��pQ�V�B*'��X
�!6�>3~!/
|�:����R|EY�&VU�$����'�ml�.ѹx���_�[���l�ص�<g�u�_ yP��"|m�cf�a�
 ��ʗW��	����X��HI���������s�%�TnE�A�4�)���8Qg�У��������V!k�T^|�A5�G���L��HJ��T��dX�]c�sx��i�Dl��hI�q���:�D�Y���ܒ� ��G?�Cmto
�1��nIA*S���\_�B42�W��n���EA܅�/�܂���Ӗ@�����K;�����~����c!���T%�ţX��]���ʝQ �[�P�2@��h;*�z.i{E�ݬ�LᆍE\C%qR�5���5�=�u�D�j�{<W�t�N$�%jK���v�����键�� �$���<�)��ۓPJ
tDbyl눫�:B���hB��E��h�O�464�ʾ�b2��9� ��j&��s��G�&�p���צ�E�f�R�B_]� O8:��9vx����&WNQߩ���g��/�А9|0��'9q4N�Ny�"�G0\�6���5�����_3(����A�/���N8
Мױ�0�L�	T'�?�q�9�:ڵ6gf��5�lr��P��u�3�?�<����ֻ�(C�tg�"�pO��Qҹ޺@9V�ϖb���^��u����&��c�N�����%l�k���-��lK�f�MEz��$����W0�����pJf�<������i�Z�%�꾣�7�;�W�
�� %:����˓C�d�<��]����P��"� -Z�T����پZ�*�!ba�<(G.GV�S�]$:�VD�X𱔉7sr$�����<\GqO�Z�^į'  
ir�g��[�0ƨ�����(���%������$�8qx��u¶�fl��2���9%�t���ȸ����3���?QF/�ߋC���kG�5�7	ϖ}��.�	N��6�?��6�[�,��v�j�(|�:`v]�$�yH?���N�Y�^�x�|bG�L�1l�(I=)`��U̠+�Տ�_����r}p��e#���(�P{5=J�+����`,���Yѩ5"Y�Ց	�r
����,t�벲��.��46��-/Q�ŝJ�4y�ò�<�&v���}��d�%��_�$��ꊨ OeS����ƕ��Q%C�����{��{M�;���|��v�ebⱺ�qT{.��!�D{�[�e֒��ū���C�ƨ���}�2��@�Wq�6�E�f��`1s ��ì�Dݳ�?�����z���L){%�X��,?��5Q[���n;�C�95d�u&!_.D=���K�;Ly�-��$��2�\CG�&7���c����9�`�����|q]�F�r7� ����r��L���<A�쓻�$a�����մҀv�S����k~r��%�X�� �ّ͟�7G
`���cf��ߜ�.LV�h{ȕ>���v̩��^�L�jvZςMi��Dl�u��9a�U��h� ��з\M�B��C��n���+S���:�H�)�IUB������̬�d�g~����~�ʀ3�$��f����ʵ�<�m~���Q�X4�ܱQk�"�+�)+�D�_�o-c}Ⱦ?��w�6�,cM��2����U�Weu\�,��"O�Ơ�N���%�D�ĸAmR�-����ڇ.'��!�4E'"����ig�������1K��xQ�>��)�?�&���*M>�*a)�qu�7�4���JN���\^�Z6�7�t���>�� �����\덮Kʋ�y���˷ �+�&=b�ٗ�f���|O���i��O�1�L�����H�v�_e$^=R̛����
�:ڍ�n�<�e@��lu�K�x��l��5�qYb��[�E��6ޏ�~l�v�_�m�Щ�s�V��!t7N�`1�b�Gj#�:�з_;HSw��#���c[J�[
��ݪ���C=SpGsX���}��<�>MA��ؔ0�j�0�չ��$D�6j<bK�Tr�e�.&2��>t��eL`��	(l��_�Z.��b��:U��$J��
I���gH�rSæ���� ["��ߤ�?���}_WY���?6T���"�|�g.)֕ ��vBÊJ��ȯ�(lJ'����E�0C��lq`��5K]�HV�i�	���D+�p��|?#mW��Z��n��r���j��$"������)�x3V�{ـӉ�
��
�-�bB/QQ���e|�����GS��EO�������t%̝��5_;N�ufD�Ed�:��%4�⛗̉N�t �M�
�2�8G��"���b�GG�)�7��3a���# &m���h�g~�sKR��x=j���-n��M�I��٣�cJ�4Ӵ�`�`-�	���y� ���7�͗O�u�&C# V�E�򃉼�Q�oA�f��嶕��bOע�;�St]���N�}5�=4�~�s��f�؋�K�ofI=��K�����=��n',J)�ô�p���3[#D��IQ��{g`���A��l�y�y#5�Q8�a�iĻJc�+� O;(�RÞ�U����<�ͻO"`�Z6�q��J���rP�i��u��K��M��r��3��JT�&7/i�7�� �odH���L�yDdF��Ws�a~�v@���,��TݳW}jR{	��m��S�á�ܥND����@Z4XB7Hv[�
Z���#����7�F
�� �F�i��i�~ѕ��B��3��SCY|�߷
�F���p�Um�>#) �=�6�E�0�P��H:��|�@K�dZ�����Bx��\ǻ�C���e��X~�Ǥ�om.�5��}'�!��z窷*�7��I�w���e�X�r�KE��CY�[HKc�4�����t�அjv/Y��S�ĠUZ=߂����K!��0��GQ���.H���q�/(���1.��ϻ3��w��/���!�� \�5%���D�����xx�e	״[�ɒm��?	=j��������?\���-\s�p�z��|~�u+�H,G\5fM�ɅZJp��° QB����H2x�N���|�[d������^����˭���?�V�#-
�V>�x��EeӖئƄ�5��4�L:y��s��>���S#�ژ���$u5����EӀ��'k����H8ۄH�:����ger٢�>R���a���{Ws��m��S��ٖ�c�#$�:��ơ}y �2�+��,��ԋ��w�dgq���L�"c_�M��4w��i����cH˂�W�d��1�������۬=�����zFr�륊�����M9=���g"�a3M�S1��c���n가�@�Mf�3pX3�Je6nk�:<h�g��K.�ֽe���8٤#Oض#$C���xb:�[F���K���Q���"�\T���c��A]�h� ���J��B���;?O��uWxq��X+�q��t��A��:�x2r�$��p��+��?��}�p�U�������d��!XD���7v�
%0�-y�nHO��A
$�{;�kc�##�;��u�aJ��+���(D�-���v"`|�g������l'T�}޻��$�%:t|B�y:O�*#W6�n���5QA`ʭ��~n=�r�D���yz�0��fj� 5�ɟ��.}���k{��0:	J�is���R�]r��o������#���FP�G�Q���$�I��3��k�Z�KS1M�������P��*5�|Ƨ���Q�~�w�u@����nR�k�0���Z��<Z��5��D��� ��Y�\����t��~V��%q �n-!�@��,���m״dKW�TG��f7��e��<n-�N7��W�e<?΂Zt���U��'��� �~e�اE������:�Cكċ�c'���Pt�US�l%���y"��a�S��`�h�D�/ۿP�t8~��$�F�<{ґC��F���TY%
nN�1�G��b�ӡ�UW���	R���pQ�~V��d�6��{��m6y�_�ַ�fڏ��	w]6�&���,��sg�O��7�A:%)tZD�.m�"��2-��M^��@c�1&�ѧ嶟�O����KT#k�Ћ<ʟ����Ɂ4�+��)��cD��.߶�M]/��.�?���v���J�t�ܚt�Ȉ��N��f|*b���gK�'� �x��{���é9ȃ�Cp�Ո.7к�φdb?�Nӝ8QgJJ ߟ��	C����]�~�Y\�����Mg˯�~��D��HD�O���̓����B�L����T�{������,�&9��'�!��[���Ng����S�-�^F�5�GY������pc<��Ŋ�'B��qͅ��k�H��p#R�gp�2\� ,�����"�XW^���5�j�CX"���Z#�o�<�p�* �:v���88z�hP�
�\2L�3�*�������P��0ɯVu�R�L�3���	"s�����֍m�;�bi�*������T��_'S����N��e��U����*q��Q�L�<2�q������{�`;�q4�ĉ2��%�f��S\�z�����:��e������
,4��u�S�<0��6�vq�b�@]q�G�9F9�K�b��	�gَZ=D�'?uZ���:E6�ݕ�O��e*q��t!t����q�e#��+�IOe��ߍb���4ȝS�8Uti(�&�vOOϢ.ȖV����ްL��S�Fk��NB�L�d�͔�/x!�"�c���h��=�6�2���--���ȥ�����[��u��,"c��Po���$M�{�:MC��,{����6S ��*p��+e5|�P� �q)���v2�d�3�1�!T^/�g*%\��m��BX_J�_[�%}��on0(���m�������ED���Z�L$IJX-�;��Qc�F�*��<�)Q�}����k�E|��~Th���8�@ �&�"ƌb�sJ�r)���eL�V�E�<���Ƿ�,6'�E�T�h��Z{v�222�
������ε�D&#�E8��r1KF~$z�����#��	WO���}���`ՓdOW*��oCc�&���/�?�.�'<��TzX\ �j2W�V���C�`��i�����n�B��QG��L�z˳�{�E�X�zT,Q�#��R�u/#�@P�v��Ȉ�z����땋�����`M�('�k��(tC#.��[�w�q�O��nF�l(:^]���m1Д�߁�O�?AX_�p	�E�:��XT�2*�F���is���g�i#�Z�'x˗ig�-{�q����>�6j ���z����,+j�L�@ϐ�6�Q�v��Y&�v#���|�_���bW�ݼ�w��/���hL���L�r�����_���k˘���f���Z@�Y��=��8T>�CԀo��Q�埫M=Bު=4D+����E��kp�Rٻ�2)a+	o�|S>���iJ���ĉ����%.�vX ���Z�*]����l����q4f�|�|1v�p��q�g���>�g�h)h��Vj���K`g`�q4bg/8an�x"Ep2}��� 6�[�L�f)B�wF:=
��o:�-�H8�8[�پ��1.�8 z��a���%�KG�ލ����M���n��F�����6CEޙ�ð1�<�? ����v�$��qK���ĉ�-u�����C�F�z�m�a�a�	���^�����.ϰ>J�h������?�V_�����?48L hc2�D��>*�1�c
n�oΨcSB��( �̗%FL�%t�0R�$��Wơ�/t��=�<���v��|��#�TW�x� ���.���[� � �w��G��K�l��35G���xm���P�ͳ۹��_\S�Ӂ��v���P��}��ƅ$�c�9��D�����`�m�}~��7*D��{|�${�ܥQ5��"��Hڮ@������+wa<D{Jͼ�-�#O��EX�̜*Z�ŇV�ט���u��j�w�)0>0�N�ij�e�u�p����H�ۥ��W��?R85��S�	�L����?
�~�l�11yY�:/��n�U��?�����э�9�T�
�,�oL����{w45L��C_*� SX}e���D�{q�q|A� �"���۷�_��!��S~�X������iPOx�b����4�YM�ۮ:���AҞ̭���/є��U0]2J �n�釉:��;>�4	�~=F�Q�̵�<�ݛ]�A8��Ḥc-�,��Ocg�,
`II:[�7�A�n��*��͕��o�#�R-���F�6�.�ޙt�y,���	�pWߗ���}� �-��\���_��3'�w���уE6�t���	L��俰@�:k�]5�{\d_/���= ��B��7資o����> KH������W�����g�'�^1�j�Ҿ���oGb��{(VY��i��]�A��Ν�Ƿ���sk����/W��h��K���-��-�LA�
���r��Φ!��v��ȁ"���7A���-�`>4�9��P��e#.���ȳr{���q>x��`{(�	7g�k���	���5�%�����B#=��${�{	��J�*`�#��c)5��I�X������t�o'�kw�>l~�u��63%��uƉUJ�֫�;���=�Zz�^Q�h]\%~{x�3.�,+���-W}L��T��K����8(�e����v�^Ȏ;[�C˯�r�!�%}�3k�(��.S�O'�����?œ�N���xv�ʊa'_k�����
[;�DN^��p(|6���G�0���}A3��#z�S��D!����5J2{��[\.�VڍNUj#V=3ڶ�����A�����Z]X��w�ڑ��\C=\WN&XF�l�C�Qu`S\�Z}Zn���5鵜�S's9��{�H�Fe��m��4����=��^Zpl7�x���tf#;���?���v���=p�gr�7�"��t��1�E��f��J���U�4<����Ƈ	k���	$��ҏ�GV* јzS�7�������q����w%Rd�؛O�u�0�_;�ƽ˪�8��N<m��o���#{�>���ڙ���\�>{�vm<�efk�q� ]���q����m �7Oa�QU5�3�iU)���`#����"{m��Ǭ��B�C��1��"�>Ag�����B/뗬uv��A��U�.���FpZ+.|~.ngh%Ғj�:��W���[�7������4pV�$����Z����v���)���#��=mbO֋�G��xv=I<*8����UH���H�-�v~X���c����0
��|����\�Q�}��m�n��).eny�w-�[���<�@����b���d�T,�X�;$v��\C��օ����A�#���r@�_M�_�����1��O7��uhh��b�9��Rtc']8/�	-��ЄR۠i�v��-H����+_hLE5<���ب�z)���G���$�� Ju���e��"��쒇��0��l�=񿓋�@X"��f� z����e�S!F?+~*ph���Wcԃ����"���n��髃ר���4n/g���L7��[ad��IL��y�G��:�z:�Q���5�N�B�� �Kp���F�/hd�K��Ӧ�[�WoН�OH��]���_G5k��R�XW��=���g�%�;��F=&ʱB+OfO'~�bs��������1*E�%ir��}��\��@�������c� KY��2O�0��mj�;q�d\J'�6C~��|{�v�Y��3G���Q<��y�<�gV��Q��oOY�&ג:H�'V9����nԱ0�70y�GG��D�����DV��e�ȃN�m���,�����s��z�k'Z�@ �{1��ǣ����59��z��r9��F���Ȼ�*W��:w2I���QU!ߛj�OK"�}�u�ׄanvB�JK�x�2�f��x�Ev`.����;��J���.��u����Z����Wp�C�����V�w���@�C�2wb҆�bª�=q�HM!��Z�~m��XX{4_���g�L���d8�$�!,)	��	��mι���<]�K{�������\*�,����
P�ʘϽWt�$*�X��AX���2>65� c�N��^U}�=�x�`L��i�;���J@�!�m#�=�z{�<I��7Z}�R�l�z��j�DY�:���!C�@K[����H0����L�mSR
Wy����j�0O*�3gI7�nJ$5��r{7���j���(6����Nm�(�s����6:ӎ�2	��9$臗�-�<��ӯ?�}ǥ	�^w�»sԤ����B���?���E�CDt+�hZb�]}����l�Z�u���5mOgJ��S����4���,��!��xi˧�/ȥÉ����HI�2�5��j�r�q��~��E�ȡ�$(;=D/��_y�ă��[R�7��j�k�L�Ǌ�1VMy.�@1[��&���՜[�1}��6Д�xQC"0� ���<Epo� m�%51؟�Any~/zKh��͙��.�wC%��n ���D� ��v��P�$�< l�T�P},�Ǚ��U/�㷵��?�=��j��iv��9].V�uј�D��*K�C��qv�%���yz�<r��\��fFj�g��H��� V� 4�_ � �p<��8|��4�J�R�u��'Kbv�h��ʅ�iJ_�|ZX�|��5ݷ=Z�C�ٵ�w�;jJ�盓僇eH}�j��@��	�Տ��P�\bH�3�/�^�$��nW'/��ؼG �"�C�`!����_����Ɛ$���R^���g|RгJ��B���Q(����Pc�қ�=�f4�}�~���\�IN�Ӽ�m	,qF6��v��^ރV�"dfr�-�|�����b��$%���N���e�t����at���z{[�f�y��i�jAU�t��Hᨙ8X����HNMg����W)*��F�__Z��6$��t7�S�#�Ţ��LV9���zL�uX�=��*�AӐ�ݮ�f3������QăHG����l�^���*&
@f�L%�܎� �`a��`����ky?d<�ϟ�Ѳk����A��D��+`j�N�8� �Ezӓ�9J&,�����))�!B�R"=t�ǐ�Kc�[ݨ�	���w6�G�$!��Y���;6���6e�i�D�CH7z�saEg�X3�_V���"p�˫,!��M��W�Mp��A�3wR��^���,�E����:}�08ӏN_&K�7���I4�+cy�ڂD���=�d���ԓ�"5m� Fz�Ȍ�����(�|�� ��&�!��|�[G�3�%ܬ��I �k~��#w;l��,�¡��!AY��z��E��s�$i����G�j�щ�)�o�����%Ɋn>�,'�׸WJ�"�rJ�igY�m����L��,VT���a;Z��ާYኋ��RϑY�|U���	���+e����KC���o�4���2���"6e�{u�q�/{�i}�ߡwO���%����'�BY���V���l�Mu��Aj<!o��5��q�.��cՆU�H�]�	�D�儵�dDl"c�׀E���̄��`�ڦ�>J�%�"�=V �3�L���f���m�.�%k���<;?��`�Æ7u��Q�*��_��2|�`*�բ��1,xpr�0n��U�)g�{a�erhE1o�"ƾ6�lI�k�G�YPG���SE�~Ħ�A���g@)�ꄇ1m�ё竩y15~���^L��cW6I���%��}hMz��1���z�z������L�t��֕�/�o[7�|L^�a�e&{lO>
\�� �"a��`j���~��9d�~]!�P�C�-؋���8��#R[#u��t�"�zF:�_��5Y�&�ks���2�B��ܝ벮7�Ǳb��d��C�~}='ឹ�����j/e,�łM*��F�Q��<�A`�)A����͙s:@�$���ыд9�V͡ll!��c������a�%�F_?r�ד_�7;"m�i�R���.��|4����ږ
�<?��h�7�"�li������[�Z�ZA@[R�w̑��6ŗ���oV,�>f/�Õ�Z����c���"��4��?�L�/"��{y/��^����6�.�T�5�PJ8���X��f��k	��}	� �FT!"�	xo#�d���3t���Y��eS�T�M�V�:���i����'�t�����d�USF*�?���w��>��z�Ň3�Ρ�&@8��h�e�"6�}�I�~��b���=����:zB�%�Iʦz�CU��F����9���nRt)��d��Z�_J	��I�ҷ�oL �51���.��(G<�·��g]Ҝ-��Y��%A�h�!H]�쨹6_6l[�g�$�G�TY���Y���#���w�6��ܗ�dI���sT9$i
�|�#�`S���]]��h��ڛ���%�=������	n�c��hF@����$��S�i"�4���3�$A��``��fPl����� .�7&���u�U��~�%�x����V�L�%��SS��S�Bj�F�ٷЁ�og�$u9��<'���b���hT�%�h,:�Z�-�IU�i&��#�T�Y��֞ L~�	ט�~:���r���8�duCe^𝞴�I�}�����Y�v��3W�~��Y�\rp�i��5Ը�\*9��y5*����J&��A�Z�-G����g6P�~���3`x�Jp4��m�<���={�g+DB��B@���z��݈,���R�1`m[�}�!:�7`{�1��V�7N�B��*��?g�oq׈���w��~�G�j}UW�[h�
a��u46�ϼux���w-
=ƻ1.��%�	*l���4����%%�;A.���-:I-�o��|R����]��Kp��l�O�fR�c����݀�k�!���5�!��$+*�1�
�iO��,e��<9;����Ě�����a5$�uA�[fZt|�On�)oxgm��!L�;�۪�K �Bc s�*���!K�S܅�!��o�-�y��UQ�	�$a)ro��I�_6�#���N�T~��Aˀ�H�!?m�O���
����>��wZ�yT���M�HtH95��z��R�9�4g�=�F�V����7R.�<k��8+֭�voW���D�]�-�/�#{��y^F�b��"�ͷ?�{V�"����Y��"�4rڤ���V�'g��JҖ̂C+��꟥-��.�-X.r�t��#�p�*U��S��@�6�k��� W~�j�N�� ����'�ACHE氮蝥�XI���y�#�(�'�Pf�����3^I��.�{g ~�/�8��O��{�a�!��8�r��1�{�����*�h�`�}���O|�F=.dz� |P�~�]}�e�Y /�Mu��(5#��>r;�� �Q�c�h��1�4�/�4g�7�>u��Y�i����;~~Tij�����J���p�8�po!�������
��F67?$�J��7�N����!�}n+%Z�èH�����iЪr"T��؇Mn9|��3�[�t?S[��"���N�J{b�9���Q�0j#�=0Fr�t����Y��m	]/��TӰ*zX=�nS[7�h�S���fI���ž�ǃ5%��v_	6��3p� t6!u:iJ��F�#|���s�VSaP�P��j%��|b�Ș
W�;h�>S ��;F�?��Q���(��s�<�w�cV�ˮ��GC�����s2�e��{�ZxX�0W-�/�b�/쨻���A����~ M������2�A�=��������@�2�G��T�~̓	t�ӫ�ݎ_>���T�6�0�F�L���֦��~������M�E�ӏ%��y1g+B�y����&v$J޽b��~֞�\4�Jh4g#s��ާ��m�W�h涑fB�����0�̽�TI��4�Ыo�m��a's�S>- ��a��r;���:&i|��۬nr���@%iE�2��%��9�J�c��2��J߃�"�F�NPM
Aw2���Fw%���v����23��}��\���&}��P����\eyE�TP�.��ʲ����m]���b�[����>Gc�+�Ku,wz�|�5��&&�rw������C�#�y_)J�s�)��e"����P��E�*M�vv�~ۨ+���5�R.s�$�2�?M���aV�z.V^��,{G�����l~v�U�ƺ�(���yχ�^��(��L!.�eH	r؟Z ���%��b5�b�S���۔���$�F��T������7���}�X�z'���:�5��P�@�����nk(�Ҥ��'�[}���#�&�"t�}���R���;�y�L�U�]+n>4�K}5~o�^q�h�8�]~��=~T���G���`2N �a��M�������X���x�e�߼��|��eʉ������)ҝ�M8�T����n�"�������+�X��1�E�������S�/�n%Uk�og�V�P�����l�i�~E�٪�_����
̰*�!e�Uԝ=/J��
g��}��!]$Y.�A}�.�.z��9�ֈ�gp�,vM��Sp���?�	/m�	4�y��M~qȂ���� �4�+̭��S%>�7Yv;��=�4��X1�C�?�Z)�%��Z�\AF]���^�G�]P����2�ׂ�{`�rA��T���ߏ��	��0�Ƒ�]�g�E'���f���dz�o�`q%�oC|`"�2�9&�Ag�~���Ki�����Wq�r�GcUl�Ȯ����O�n �� �d��p��u8"�8 �@:�N�A�yъe���X�%]�`��XW2VE��b���FF�^OEq'���&�(9o���ף=W�$m��:�%���v-Iz��7�8J��̇!+��['�Q�5��F��]���qFg����4#S�d~�&/'�o��|K�eZ��\��#��j���}�V�x�A�	�Lk����9L�O����4�חo�"N��3MT�.*�i1�i��6B���VLi�?�����9?���>Y��d	 8�	>�cj�.Ş崍���>�@ n��)�Ei�՜���5ـF,i9��(��y�I�[����S��j�����!��̮w�䲶�oVƍ/y�h��6or����Ș�"��+U�/����0��O�e˿�C�!���~
?��-��Ɩ�h7'3qG�}ћ�k���PS0�A�7��=`�_����(:���.]�h�oT�z�9 �7��T0v2)��ΐ�P����%���a��]�ť��Aa������$�s'�Y8Y�־��69��s^��'�D�fn��i	��Un�x���~��u������pN���2� ldAU�0��7�'�kE�[��
����5�uR�ςW-Fz��Cc��2tI������fC1��eѬ��\q��R����L��� ����q�|<�oz�zNW�O�)w���p��ӽ���並Μ��˵�V���E;��sq)�w��k�h ��!�B�O�	�@��5�떎3�䡶4��Nɓ�$nG������ho�O��Rx�òF̓��M�8���B�&#_�eD-Ĉ�$��-mg�k���aП�׬ ��a�������Fy\MV�.��R�c��?dy�o
Y(���6��WSzH>��&�
e��T����7|�����:��J�	�c��
r�!SY�c�)�NB�Gt�aqG�8����_?AKvU����J�J���
���a�+\1��l�:���6O�Q�hf9dX�~2
ԇ�m6�B󘞉�HR��B�<��D���}]y�YV��F�2^���z�;H�Ĳ��ߵz�4����W�ǹλ�%�&N�-��/��2Ńm��[�J��ךkʉ8#����%3q�4��y	H8�2i&��W�))�_Pd1��Ƽ&�mI��ox��;>?�;s=�Iy�ӹ��%x���4�4��I�\���%��Dz�A�i����πP��;�b������*W���S�,��&��
M����W�����z�#��o�½�G���5�{z
Zy0��pK���>�'#e�e�Cyj�K<��R0(��ԕZ���O�3��(�����#��'�V�����
:�S���w}F.{�����
�Αj���1�ѭ�m���?'$Y%5AjGĭ|%�(�(Hib��;pew&�I��,Ox��g1�Z�^˒����ɃP�f�������B>_Bh�;��H!�[p���X����%��9a_���wi,�o�6�ż�H׿p{����^����v�*��.�����u�*�op�0��C��c��F�P��:�3����I�z�����[�<V��	�Ґ1�n��j�B��8ӱ���\ �t�=@��a�ʭ�FKx�QI�F���-(+Ì�Z��X�Ĺ<P9q@��E�I�Z�Еƻ-jײ�G���}#1��-[�݆������I�h{��a�������r�1�ܘ��֨	q�{I�~P�X,Ɨۖ,%�kz�,�L7���!���y=-'�P	��(�Z̊b� ؑ����$yF/��!���Y��-���U���+�Mu�,oK%;��<U=B��"NL���py�K���jb����fQ���h��Г����~=�>��<���N��]�=J�� )˲��A���A��������̺A2�p�"�hJ&FpͰ�=�u��^C�vM���!��i
η�� ���#~�$�Ŧ���i�H#6�������0G�_D*�����υB'�[Qs]%Åplʉf���7���W�*#���n�7�{��[6r=����R�O��W�8�F+څ*���khA[�#�Ն�ſ/S׺���,'ઑa�v��};o��l��p���MG_!Jӕ��0� 
9�^�ܥ���� OJ'F8���Ĳ����q�жa���vMÛ�ȮD(��;j3��)K�%.��K���u�4+ϵ^9�U3x�g��UQ���=ɹF��qE�?Ƈ���-�������K�B�׿�A�1�	L�>^�S!HJ�*�q�G�v�e��L�I�����Ds�ˑ���A����l�:���߀R�'���X���Qt�b�;賯���3;��F�ͤ�x���Y�I5���O�%�K�&� '����;��Ig�l�!ι��'ۿ\�E�t�]�i���aV������O[�
��a�B%?F&�nї�N��xX�t=���1�|��e@�Z�����/�A�(�`�sV�2%Uٗ����'Q�Ho�ڛ� r|��.}Cz��]��Z$&�}q�M�!�� ?qq�(<�[,�lK�(Mn���4�J�U	���kKs�Lp y}v�P�a��:�U�χZ�6�+���l@������W�W�a4f\۸\q�I��g����Xa����"^�ɴ#�D�����դ���d��QOqj�+v��h�~���T7�:#g{�_ƞ��_W�0���^�X����o߾�X�Z˸� =E(�k�����-"���a��Z;�M�]`�Y��}S���� p��y��2�,�o�V~00��^���	�S�w&��qR4	`-�O���^�]1��v���w�4�6�0�����'Ѷ8)�e&�}#�2����i&������R�ZV~RRN�� ��_�{KZA:;���x~��puC�y�1+�S��� ����Z��u��^Vl�؆{f�ҫo޳<����J���#?����+�W���P���w.�)Qu�����5B��$,����6<�f+̍N5W���%������f�����_��"Q?;�ĺ!��}"9��6�g�"��G�����#��`�����tu���Ћ�R���k*�1h��~:
�δ�n��Х�aє1WFG�{<AW�!H��8ҿ�͚)/*��σ�B\<����~��&	ۯ�ÿ��2���)�Y8B�c�W���N���-:�	�� ��A�'b��l��|kn��8~���Wv�ʗ�\�4|�!X|b��$��B{�%�v�	h�18� 0h�.����)6�Ȣ�+2��S��E�ۀ¦��x�wH*]�&��m:��>�Bm���\#\̓��/L�y@��ZV�8�޶¹����dc�`.��4�U�q���i���F��N+��� ������u�;�,��c��Ff���K17�%M*�G��-�*`R�㐧'+5 �n��?Z��Xl�M<�J�J��g��:
�%/��>��2뼮pV@�����%�b�UQV� �ۃ�N?1��Hyp�[}7�̤�Ʒf(b&Іk�P��P�gS� o������F9
�w�D�u`8����U�6;�l)�S���T���;���>�z��nw�X�D[����8`d�h��F�q[�6d/ă+��I����&�DbF)f�_~�lI��y�bf ��g!�Ki?��`���6OQr5;�_� �Iч��iLi��X��$��hĮ��۽�RR���i+�s̄�X�FFus��㮮�
hq	�P=n���̉5����E������z�n�W(�vA�ϸ��U���7	�A�<�Fk��O��p#�~u,�NJ;�<���4�\U��t蛄8�S�X�(j��%�l�vw���A*��dOp�`�9?c��f�$��e�D2�#;����N�Ѻ3C���h�K0!ҙ3���+%��~c��`d�'���n����!�����������(z�҈�ݍ�D�:DL������q�1_��W���t�z�*���٫o4|Rt�O3��2尬X����b�^�4A$*��
e.�}�i�dl�)��	���e+jv�"ƄMj����5
-gZ�Y2i�J�A���KW���9���b���q��v�U����&�,ZfST� <�KI����K.Vts�����liPym���{U���F����(J�ι�|�!�/�a ���I�O��zMz���kYX{̚�E{�y&�������jm���	^mC�=<�����;���հ���_ڔ��b�q��e�K��5�Ι��'��fuv"�d��>vq���)�y��Qz�́�β���~���E�9����=t����I���W[�HB\��zp<��Th��˻��G�2ț�X	�� 8�ԝ�w3B�}Q��f��*��o�)2��Ik��l[�#Va�C���pm��Oׅ7)@v�w���4w�\?��:����Ŀ>�㻎��
4���?��)�q���/�[����CG��y§�8��P��8șq1�>G.0 5��È�ݎ C��7�2w�b�����o'��T_{z���EЄx[]��p�QY���� !p�������I1��f���OE��OȜ����wY�6��%�y�ߜ:��7s�&�{!���)���4��Y(��1"�(*���f��VA�UU�L��Y��v+IT�럈�f68��7!���p��9�'|)��9�WO_& ��Z���=*=�V���ZZH���!,:��[9��UF�l&|�9Orǵ�������������Ia���`Ս�z2�j� :��!Z�R"��r���1�SL�gl�ST���}U�ӷ/| �V������t�"������K��'���d�(.���^�u�K�d��X�������s"�w>f�Κ#�v�V�-N)\���������u5`�U���'��5����59ڹ��	Q�.�ƃ�����N�<��C�-�Qs�hc��F3��I.\y{ǧSI7��3e��O���d�7˔Oy7o=Ŋ�H���`���oH�
�)-����{��S���Ai�W��^ī��~K��<aHo� ��=r�L-����7�W+��N4�}�'ԋ�JM�3�"lk۫
��}F��x�/���H��i�m>��%r6J�{��]�$1����ΰ�ĬN������AI�L������G���M\K�tj�����g���59>T���,Q
<�D������E��4%��]W�'�GѠ���`�4s�u��S���ј����y�W�������j��˦x���j_�������~k+v��)�^R}K��Y�������wV�D���uaXI/C!a��җp�P�_��z�z����K��9�O_�5��85M��/�׃��i��E+N!�6Jy��Dm\���R Z[T:��TM�y$m���,M�n�9R��F�\}<#�8��ba��O�����xt��~�a��<��k����]Ic��J�d۽�݈�n�<|Nuq�����|�'8)q܏4Q(�����3	�~��0��E� ���Us�B';�3h��D�F�0�PE�pi�3x<O��r�r�ݢa1�&�1��P�N�Ba�W�@�kS��/��|�M��p�$�fs����n��oc[���ߤ)�$K��g�P�	��i/��/�m"{����\d�y�����?]���}�87*�C���e����a׿��
�9���=i '�m�NjL��y�7]u���M�`��h� ;ZDӼv��h8UN`�r$�^,�~�p��w���4�ú`2B9��}�R-O���,^5-pi��{�z?(bɯ��A���p�@n�T>!{�<1�(�-+l�룠5��)M�	�.v�O�fѩV�Oqp3G�� k�.��&Cp�Z֎]uB�`}�1���yJe�N/��ެ����Þ�|��D�\F�
�i1s���>7v����j�)�]���_i9'�W1lf!m�1~��l���	��8��=�D;���|�y�t|Ƣ�>;����M�)kNSU��"�X���I*��P��(��R؍x���m{(*
LΑŤ:m�^yjj#�]aZ�T�,(Z2�4�� k�$n(
zD����Wn���~׻��� �g_.���6�{:�r�����x��vG�>�4�Wț ���>�v�L�:s�_���S~���g�0O�~<H�r�7��ruw��6ɴ ���q����*-�ͧ>�6 �M�����M?�G&T�u�B�1�X��=��..�f�s��d����w�"hH�Ji|������N�)���Lv���GP�62�H��1a��X��v~5|�{�x #�;."��M��uT�y�u��<��l�t��03���¸��q����L��������7#���Ef���q'�7�p��������}�rf�|�c�q>3��α�]�<2�+�m�L#��/�F�z�o�����v�cח�^�D�s0^�IF��E�Мa�0�ܿWa��+d�g�������\�����"���
�C�bJ;��S_���v�.s�-���i��-v(�J�T�g��d�dB�Bu�@\�Ƚ��g�oWls��HO	�_<�O��
ob�f��8-����d<�F�{�B�ƷP&OeO	�!��彌Dg��U�pn�֐�p��j��CLa�K쨾Q؃�{���<��▌��j��x!*�2ʜ�p���Ɇ�h��qѢ��f��#�#N�>�;d��R��r<}�m6�%��/�(if�iƶA�QZ�
�����	���H�c�g<h���D{u�4�I�F\�y?Nڡi�<��֤��]���+����sT����:�9�Z4���[F�S@��΂<LO�0�>�}�������3�/ނ:$7p����W�x��8��l����:�cA�Q"z7#Y�w��j�|�ຄ��pr�O�a_Q�Jꋉi�R}n�M;->Խ��W�8��]���.�P�[�݄�љh�[����D=��ć���iG<�,
ؚ�Y����a���42lu��iY�n��$�ՓO�bF����נ�p�ӕ��l�(ir��5g����;V�1�q������,b���y��Ϋ���*�%��2��$�����r�#2d|�)֜T���ⷠ<3����ԵHx���?�C�w�m�X(�p�Gw�y3(%�"�i���6`d���xq?����#�b��d���7���T+�;1g�	��3y� +i֢�T��|��/
���ܖ)2�P��������� �W�հ!Voĥ�s�6;�$�v�g�L�x�fܘw\஖�����h��c���[7���ـ]�C�hg��ӊL/]L���������+�<N��fD�'�E�?Ԗ�� �]z����1� �q���_u�KG�TyK��67;j-�;��]P�f�f%��v�8-��#�9��G�Gװp���Z����OY��v\�SQ�E��[QϤu�7�@	��)�O�!�{
$E�$'>�}�
���I��t��}�pAߪ�����u��A�,�}�ňq�e��p�fz7���R�o酪�'n1��������L��	fp����|�ƃ�� Ǡ��	H1ネ$O��{i-/a��Bm��J�%��K�1��*�+��G�4Fm���Š�Z��̲� �I��2�X�s� �����g�<��6k��:{�Y�L'�!�ss+5���OꙠ�MC������̹��l�vq"���m��z���P-ϦvZ�[�ᕊ @���W��qi�߃����	��J�g�g�M/
pU�,�?5�RL��02��B��Y�2�*U3E���G����X8�6�(����O��ꤟ�c½Q#��p� �O�q�`;�sD���J��tTKD����>�xb
�����'f@�dmJ�e�h����m[	�S�.�w�eF�ZU{~c�1��Z��~-���	^���U&���s�V�z0��3�bUg[�\*�r| Ƅr �1$1����r}?Qr�1�q�k����CL�t�I'�������N3�K�!��WW�󑫁U��S�_%�����g��έ�w����A&�δ�"�����Y5~���/Ps[j��i?���Gt�j@'��%o�+�v|rf�f2��[#<n��et�!��|�^�C.�>H�(�+���-��D�*k��P���o/?�<����?u���ε�:���=��Ҩw-�]��|e�4���g�>��\J�|��d'����e{I�c�y�Zn�V�*�X�)��ѷ�Qn�*$�28��f�&�B\�2v��?r�H$C����uG+���������k��1^ �4�o��a�&���^I��Dm^�4mf1˪��F0w>3�kp���{w�l��9�`�w-ٵ:����CgX^Ǯ�?�k�B"T�.%���|�����Q-�&(M%�',�[�,5о܉R��G��,�<�ܹϣ����ME���b�%�	�Ŧ��ź4��5�NPbWX�@D2�/{&�$�Z'q@>�v`I����֖°3#�
ǯO��M��Z�M��)�æ��3�xR���Ӟ��S0�^��_�Z��b�j $T
V��U+���Y������-LRڴ�f,V�阮��#��4�U��P�2p�F��	���ISSɧ<�o�����Uј8�*�%�Ϯ����Q��P��',��f������3H�U�ǕÉILx[����z"@�a-0��,x��t�6�������uQ�6 �s���i���;nl��o�7���� ž΋�Us�AZA$�DǄ#	�[,���uv����+a���7.N��S;� ?��
Ͽ̢����]'�B�((�X,����PG���t��S�8r3>g���~�$� ��۔�I��iA�H����l���˛��S��%�7uL�8�M/[xӲ�#z�� �ZN%CKc�lݹ'd��+�i?A"�E�m(
�*���P���c��8]8�����e	BXzWv��`�Θf�kq�H5O=���,�C�{Á���4ˍ҃YÀ>KX
��gǯt��H�K��Q�"o��W|vcm��J�	�����Y-�%�W~��[*
���{X�	n~��� �v=E�ߐK����s`���{���Da5�aS��9g\���	�$��׳���/h-��۔(��	u`y�A;�y��핻M8d�ـ2�z�`V�NG��(� o.�Ț�	�!ٔ�5���B��t-�i���[��򇖅��IP�|��ᰧ�ei�)�XI�@���qɐa�xz��ܐ}�}#��]Z����2i�:�`�C�.�$�T��n�%�|T�Q��g��F���G�=�>u�]�f��7�+W_=����О��,�����9��f_�L�Ӗ�rc�F���xes�֥O��!fv�X
9�1 �m*�
hrV����C�?dՐ
w+���l/v��7�̇��!�ۉ`�e��f�Z�B����%/�UCud(�[�����Ʉc�����?��K���~��z�p�0K|����p~hTܘ,j����ڂ�,���i�J�$���f N��'���04���>S��Sk��Z�������Sz܇�F�v96��0+"z9��CQ�A��T�%Ȉ�	�H��D��G�2fg�xkU�������3��" �Ո����7��-����;���H?����[�^�J��� �Q��c�C+��H�t�v�A=��R��{Q,ߡ��#-�&��4:�~�������F�!\��>)<��$g5y�jV��b1�.Q�4��;�
�.ظs,�nҡ8թ+ťΆ�?ퟓ�>��Zx��ѿ�����mR�&�ʚ"�˝��E~@:�WvI�����Xla���7��Ǔ9��(���eJ�MZ��f�z�[=������EI��P�y`..� �e��K\�t�_��3}���ې)i4(�d��Sg���WҚ���=�IS�D��~�,<߃��O��q.By�,:,9h]�Y6N�@�`{��2��F�����M��09_��Et0 ��б�|�e��&m���/��DM�1���'�k�-��7zD���2}��N-L��a�pr�8ғ3]7Kj��A�RyV��*�d�M��;Js����|V�.H�5��������4�'a�j|��r�K�.�E׭dϒczU���@r�cERd�o3��b[@hذ��B�@�-�A�O�hQ,%/hzB`N&nm�:�oy�_�&�����r(h�m]���x�	�"�m�T҉\��Ѿ���b�0,�ֈ�i�W:���s>;����.��_��6 N�@�X�2��S�.Įr&���Bl΂�T��W�}�e�k��ͼ~v!d�
	�kލ��YI�%�03U8gU�{�<^��X�H���.���	�S��C�@@W֗k��{�]<�m\�JR��/Fr`� ~� 7ĩ��Sqr�tYMu��P�3��m�J;EU/��S��L:���[#�_���@5m4�����I\���������G_��;#X��yo��l�[9Z�B��xB=�ܢ(����,J}�D�l��IۡV�co>�+��t�8�LR��"J�+����	q�łcՙjX�M�*dPW�� ��(�ڤ���ACijpR��7������� �H��ow��܎�3]zӲ2�b�ۨu?�ݭ�<�/p�*�s���A�*�a�S�Ͷ�ׂCT6��K��Zis�@%+�v�W�c��,94��V̱ʃ)��Ep2�Gz����ϓ`��+�T�|Vb�!��B��^5n��S�����m< rIs�JhY�8NϛRJX�S��K��H(�t�Is:2cj+�q�� ��haK����کF�H�a 0%-�oѳȢ�!��u�?��o�p�fv��k��|�s������6C��o�^����d4R���-��f\��Qu�i��z�L���+'Q
�v	,��l����-mǳ�J��K��SOzs��t�T��h
*}1fR�~U��,FX�V>��*��`%��.Wp��&*D5�eE3,�	�S�!�˓�s�DQ�e'�foƇU�fa	�a�ٮ�w��ġ�iYQ�i�̛���*��+�b��7�z�/���o�Ǔ�xOlC�b>�z%Nh�aZ)<7�!��eU����HNV���Sn�9������s��|T�#̲`.D652�Y�p�X7\�-�G�З`	��K�Abd�1v6�KZ0�?2+��m'��-�Ώ��1%HN-
�l_N2�`T0�aR��7��lQ0D��|�#L��D�U� 
]�|�����<rw�� ��\;T+��l��rm��V��Bb��C����ov�[Mu��r.q�'�'�Y�H=�n�����G������?m5��zAO�V1�>KP_�g
%i�Ï�����ll��gP9,<gQ~�n���)/O�S�@�o�sW���4��D?	��M�ZR��u��%R9�!h�Z�=�\u�J?I�&�Z�W��Ip��7��yt�J��o�|��|�%��ejF}��]x�C�0��	�N��S3
��͋H�L�>�rc���˕\b1Y��<����+Y�-�ʆ��v-�B`�ڈ�[3��V��BJ�t�����f�J��h���%���A8�â�K� DR� 1��iJ^���Q�dPL�^�@ �X�+i�>�GLI���}I.�ip��p�cr�u�k�����X�_�ό�Ltc+�ʶ훢29Y��(@��E5��ҧ�GY��:�}�9Կ����� )�:O8�����8�'�Z�bэ�Ui�H��aj��!)��AB�^�l���S����n� �J�r��+�:-L�뱨��}��Ch�K�s,`�tA���_do��p��V���<�?|��յǣ�ȟ������K���u�^���_��6�	ŝ%������9KD(��i����1��$��s���P7�d�����Mu��DL]���h��![�����>��J�1f�z�4 �����=��vl���Fk��s%�z����Eʷ�ҽ��9&Io���6�G�k^��ې���.Z�����t^c�����R']��C�|(��6����eL�9��s�h�PC]�H!��*'���v(��DL������+�dGu�x�N��`��k:���AG�YF&�A���-�����kTJi��ܫ/�S=\��RߟpZ�Oq1�V���C���8�E�^�G&ַ��l�,=��?�9y_���I*��;����#)�+/�\��2g���k�1�A���V��Й��p���j��)y�Z�k`S����D�g�y��Z�X4Y2��F\�z��oVDL 00��	�&P�N#�p���-b`�&O�����U�6O�ԉ=�"���ŭ���
;L"� V#�6AS:�np)��*i9U�kJ�N�	��z� ��?Nr��V���-��+H�+�z��O���U�Y@ۖ�t�����?@�F��S�~�~8��L_��֖��gډ�7�4�)���%��@��f���²����s|t6\�lꁫx�c�W���Q�*���:#�y�M`���ަ6E`6�P4[��/Ʃ�,�D������ڃD̦Ac��T�|\���`0�s�).���P�	m����FƣX��=�p�Cǰ�w�5l�� �:�L��E#�N�H���ܫ.�����5��dl��]S�v�,k�*G��{Z���
L�O�
<A٪��o��ƣ��d���Ģ#2=�Mo��YE[<-B*��:��~�:	G�{�����E�dG��bI�j���A��H)�r�8B�Z�T|��g��h�F!���ƣ7{`��.���|�39X�~��9�mD�1z-'$*)�Nǁz�>����F����@��a�)
6YNk/��9���/����5�Pf�mt|fIKߌR��j��ӝ�-׍�y�dY�#!�)}^��� 
�V�(�O��i3���2�o�~���j��Oh-�����r�0h���^�#q{!���E�M�N���s��G�
��������\��)]���9����rd�T��O�yہ[b,�e���? �o�驪]Wڦr��Ͽ��4-V��sʞ��ս_��3��+�5J���Y�&������B���Z��Ha���)���ך����,=Ծ�fb�"��F�K�`���#s�����4��Q�'��d�#���]�h�3�$����J�<�}A~�V��J����J���o��㵡_��ޤDQ:��,V~�Z5�"�!������U��)C�X�5�y�,��T���%ޘmؕ72�t�l�Ո�&�>�O֣�h �W(Rl�Zrx���7��^ɫ]ʆ��,��79��y�1��<5NшrjB�K����q
�@PN��+Dq�%�Ոn��sJ;�vfٽؕ�M,���Z�[�AaK���7n���ۛ!9?�|������h���uw����y�{��m�w�ٕKL�`�ڤ��|m7uU'v5 �xl�"����R0�`;=O=�!��Î�n��<�GG��-Pwv0Lv�5��"��ͪ#�#���P�22�38����U�a� �Q�UآG���/ ���'�����S&��Q�XG�5��J��g�.j-����(4�Wi�lfs�Go�/�P{[�����Im��M���g���6o�T}�wl���]��Y��$���K�!��+|�������-�M�������2`[l2ھ)��x&
���+�v��F1�AD�x�(�s�_�u`=M��� ���ueR������[np�YH�(f�X�[}Ʃ�0�����3���H]��ϒ�Ԓ�c~�k:ނ8�������=�� Z��,��C�Ya#�p�����LT0Y�g����� ���b����;�V���#T�2��Վ�������͖R#����]����y�vx	1eM�(�ɉ�d.�L��f*���s���z�肪"�������+��c�1�IWcr��p܏$`L
��?�P�==���v��T1i�Z�*��d�e�~���"�q��󁞆��?o�ō~zu ��S��X��~�_r���<�e|BR�pmr`A��j�����U��2?�TP?��U����U��wyC|�>�߶-4B�&y��
g�"�S�ۢ�/��r.�!9���4�ƇmfN*,(���l���o����F_J��jðP%��&��1Z;��}B���`��A��Ф��StY3����
�E?����������(��b  n}$�=�c���YG�y�Z�t���&ؔHO{��y�0�m}ƹ��~�^7*��s�� ��/;��E7�4R]r`BT-m�{������ڤ��"�S��.L2�X��꩷S�[�<�w���h����� 6��oD,k���O�喴7G��QѾ
+kl�S�=kC�O����Y�ݬl�]�n�=�p��3��;U=�oi��� ���i4F��Z�����o�J!�lΜW�=j��mA�V��]Bܷ�T�NŶъ�t�G��8��f����D��o�HDBS�>Ȕ��6����ؿh��U��k��*e�\�sX#�g�ȋI��l/��;h�����y�z��;�F�&�pl�v>S/�9e{���Zx���Pm��>���,B�I}]�������%uie�F���^���E�Иs���{��c�mQ�_���> �G�j�}�%s|<]y�"�~ߊA|�r�.�X�l-�<@��e[-8�F�\��toB�{�X�7bY������X��+�e �1�]N�튨AyBz@���R�!Bv���)�g���~��s�v>F9��gmh>�ߤ��\a`�~g�#��S��؉���r�5���7J�2'w�j�'���lt�+���F&��oڈ��_�c�֣��Ȝ������x|� D�[s���	.:�c��p�M�0_aK�r��e�c] z�3<���eyH}��%e���G��1���~�z&��_�VԒSă2�� ^��ғQ��Ts8���s����ia��PfmR�0w�-_&�>�D��'q؍��(�����z#�/�?�v���"P���/$++�o�<�*Q  �������@���o1
$��.zR�AZ��ӕοd�_�I�QD�!X��\�Ϧ�nܵ��Hex������`�Z�޺�W��cca ��$�� ��� ���w�)X����6�3*��:�7�$��)ASLO��ް�Ҿ�A۝���/E{z��ɔʣ��!ޏG�t�,�/W���:�H`�H VD̍fI�G8J��m6(����̛����y>17���ܵT��ڏI�l)��חh0�ZE���(,�d�����r(D�o�f���$�p�����fbBͫ�Wpel'�8�B�nR��P+ac�xD���A���pe�wWk��&�J��mF�_ƺy�IH�3�WK�=��\�H��X�/�;��g��܍:w������b<�M�(c)6
��}�N(4���̆��ب�]�n�KD2�
v� ��?xrD�n��Wa��~ ��-0�j�`������b���մ̳r�������P��v���ފ���0m	Y����n%�E�E�ފ�U��������+�G˺U��;�q�VF�N`B`1��o�M ��Y�GI�ȑz"�-���W	���s2�V���J��E,\K}�Mw�����z@2�O3g���kI��V�W'�+^v�"���ݭ�2��O��E��N����1q43�e��?�s.��[�{���Â=W�~4{&���n�	��rT�~�h/]Vv%}�<E�j��+t�{�C|�kԵ�Ύ,�����2�n-]	"�|��J ��w^P�Sv�,�%Zl�e�˔��(v����0�Z�ABH�T���TE�d�ȣ���!��`��.�R��`⭱F�\w�N3u����%�<W�% ќH��"ZC�.kA'���$�4&G���!�Q�)\�^XK�(�5
G��AU�'Z�o�} $-2��[�i�s�7~\]�/�_T�}����_�N���a��5(��~�e���Jh��M9)eO��D��Y�$$�Ȟ��0x�/b��5�XRy�s<d�P/<I�3�\����[����&}z:2C��}x�,�2���e1> P;��޽p i��׶���e�r���YjM! ��k��ǅ?�(����vݶT�$�Q�Ul[�z�=P��ebʚ�3#[.Y��r�Y'�;��b_��y#�� v��&o�:�0���{y���B�<�x� ���'r����WH�&�4��A�F�?c\\5�Q���*��e_�um�=����w?���-����-�s�'Γ�1m qw�Šc�	@zC|�K,����Qh�mÝ�s7�Q[ݻ��$��c�SF��p��Yy^������hO�O������$dfY�s�Y�K}x��Xv5��j<����(�6�c��:�ިQ\ܚ���(�|�S^�ߤ=�IS��b��4J_bu�@���Ѱ��N2
���'^#���4�e�<��?��hxu�e ��B���}�<�BK㗺��MN��3.m6��fP��w�>Zu\���g��T��r�J���+��E%�=ڊ$'f͋�R��K�n��\G�0���N�/�9b�c.`��?�䵥a��9�zƕvɯ��O?C��Ҧ1C��9��2B�x~[c�`��K:�h!�a9�ʳ��f	�QX/��ȡ��0h<����"K/�A)��ؖ��t��#�m]����b���
S�OR׺j�E�J'���/I;h�����b
�WϙB��pj1*t䃬k|h�&��q��(��G�����Wsoб=�%.�lS,(�vt<�q�-�qwf߯Z�Bܟ�'�PB3������g��5�+ >Ԡ�W��*GJ�ZfpJ1L�AO�k��Ƥ�V��k|���Pvt�]d#-U��؄��,E<YS�R��
�3�m)~�=øQڐ��j�_�Qt/�Ji�����| �`�z��A�W6�R.���I���uZ�ː}��Z9�xY0�����1�p���p�3��9���_�C�"��4�`�@$��@ic&�g5�ꎈ�
q�ZT� {xv���$�#|2u��
���
;t��g�N�xր;���~Іm�U4��0FhXU-�	���Lx�����J��'Ѯ�R���$hz%:(P���>��4�3z�(�N���׉0��jVU0o�ԉ>��o�Ð��ێ�i�Ã�����v��t�D>t�$D�L�+�|u��G1Pzs���K��2a���u9��xH����y�y�)�m�腎���ɕ�.�T��*�zЪ}�׼RA+�ƽ��a9�L�W��	���G�`V?[e������ʠc��1�¤iBx���r92b�,�Y��Q=��uO~kH�1p<�]���9¦����+�0���rՔ7�|B��N���:i�QB�;EW�_����Q�
v�kdo��PЀ�9̐b?�6]�"P��.k���������.����������/��-�8���c�*j���gت�Z�����1z�a���V�$^���3��\
��,5-�:�d��S
���x�P*�\�w�FqZ��K����>��/�%o������Ǭ�'�WAޅ�Qgn��!�4�f��Г���ӥ���W	�{�$�c{s���B
U޸�{-ة>��8��*Z��xm���^�N�@�2h1�/��С^��^�+��Q���@���ŝY�~�����橪�����Jj%zp3.Z[+�MT8�_�YC��4j���.X/^ғ�i�CI|��9��-����*��`�����+p#�PwY:�t�:��wQ�H���оn/K��c���%u���s�}n,|��R��w����2�/�T5}Eвa�y\R}8�ۑrR/gt�(@����l�L�I#۱��c/I��D����a w(XZ�րRN���[s�3�0��ìDڣuX�)�x���@��q������C���EI�����N؁���1^E�	>��`�����`�S��H�+h��<o# �JI���,�(<�
��`��cA��f�Y���)8 �F���s�H%�`�����"e�4�}�F4��0�)����C�+����txm���ޮ��N'd]hd�j4�&o���Z��I��7�M�*1��x��cKrUDjdN�F���%/�\N�3��)��4���Q89lK�Y�eF�0���t�����$�C��ģ�/����2��~Ia�1�2 �)b:�y@#�/�FqU�} f����@���l�)]3w^��ǥ0�U��.���*D��i����ۯ�M U�jO���3m���5#��W�9:�'��:��̣��ך/T/�y���i���5�ݞfO����������a�_h�����I��+N1#��Ґ�6�
-mK�{��hy�*ߛ���C�CJ��o.�B���z ���7�D�@���m_��$�<�X�DMX.��V<~6�-��X+8@ �G("h�Q3�Byv��Tj��Q�����)��!��$8+��}��
z���?�[�8r ���s�>{@v����$Dƕ�.�4k5�bp�����,Ս(�%��xvX��D"����AѺn��a��lyK��E�k��,��Ϧhl�#b���$��7�xSJ�'���q?��5iz��%<
���c�n�gͧ�Q-��|~���z��<s�����!|�\�R���앉4���H�Ԍ4��J#�Y0��t�d�@�T�g�}�{�f3��^_�{~��'so<�L.��{/C���+Tc��9><��.��I su�t�z,�������-q�k�ʂƢ6���X����$�??���"0�8iԼa7�yz���>~Q��@�ְ�-I�!�/�_��wJ��*D`[�q鿸�9G�QpSX�0�(���d�q�ly�Pڂ�ϸ��DX�� ���Է���(S�:a����T��o�0p�B�ã��%�F!�3��Xٓ�E��T����0��Y���If`*�
�5�-��Ա��>`�P�����#�H�H�N��f�f��N��\�H@�dF�Nx��	3�ky^>Y�.��Fch_�s �q��+��������V��c����<�nX^��mBA���
�*���Ϭ8���?Pi���!���ܥm��*���d)�,u'�T��)>��I�Od��MP��Rs$�q�p��*���V��d�y��z��58���C.��sM��������fʠ�X{��O�������3n�$X�����j@��DM�'1L�7�1�zZ~J �w�3�`����l
�ۛCA@ID�5���#��g�<+����u��[���^��q�G/`x@�N�6g�1����o�h@���'��O����i,����~�h�6Ґ���-�2`#���ɣV�l����u�$���ƽ�</�wQgc��OV�˲r�e?:�w$�O;�w��	�鎞���d��&^/���Vԥ@?iZ���=���Bw�K۫���T,��'��~�s��M̔:�J�� �Hj��a�������g]n�pf?��	�կ��!χ�lDXq�NH�p"�Jȓ�&�������L��^�F���mM�`Vs����&�$n�}�0�5%�-�ً8B�
��\>��yz�>�t+YՉ%�2S#��a�}��U��x�Y�n������Dŋ�#~OI;��2��9�t^Wu��gO�&1��Jj�h�0tO����sP��^��J�Y�}V��c����:�Xg����a��e�s(��[1w�=fd�Ǹ���0�u�G�wm�:l)�;��=�$͇k���f8m�~�.���F#��Q�N�O����"5��*�Q�YbY��\$fE��(��+�q�{Cİ��0�t �L:uޞ�#��Hk�B/j�-�$�wƏ4���E�667� ���x��$�r�2�Y�X�Ɏ�"����:��R3H|�o�ʠطXƎÞ#���{�UQ�(�n���K꾜>�UV��2`s�F�_���]#��� �y5]1�gY�RX�+Z��X�`?�+�Xա��K��w��
A���h����8Q�G��:�=AteI2�	d����r�x�>�o�2#C� �I�i��/$rjbr��N��KsA�+2�fރŝp��L�בM\��`�/�=֣7�u��gG�k�
U��ܚ+p�J�p;��/�mC}�f�&�؍�@EhK�C_��-��D�lyM/�u�&��^�J�1��Y��a�Y*�<��
�6tuext��n��� �ۇ, �8��;fp��8};�c��˱3�K�D�+��B!��{�[�7 r���fR�5��6�m�[s���g~��"�	�c��!b5*Y��N�W�ߟQ�?-}�C�N*�!v#�o����z���;s_"�W���Z3Y���x����k���촤/�Iu�V�A'�U�v�e�2��Q_�,|��0��щ��[�;��G�P9�:y�<���3,:��g���L-��/�����A���۲} ��|a6w�,�DwaW1�J�ѯ�J9z�k�:��b�߷���w.4Uh�	�ܡ�R���0����Z�d��s�0�A�z�i|Y���g3�I�R�N�3Dw�����-³��s��1����w������	ANjQNw6l�:,�R��������$�i�=�/���t�8{v��ov8��:�G8�y�X�J��g��pI&)]-�R�;r�$�U�>"zJ&d�4���y͛_,)Y��⇑��. 7Lӌܓ��n§��MaGTTf9�_�sjK�idM�K[0�����S����)�t����Z?d�4�\�G~P=Vf1����
�JsN ��:&�y�_	}��%G���{�F�fe|A�,r�p��Ί��:J�����Y<�,z�P�t謘a�Ul=tXFם?�Z�F�F�PX����(�A^J;x^fוU��Qw������o:��*<l~�TǞ�/s�`���G���0&"[��("q�N�\��`������8 ) \ӟ�Em{��0��F��\Ӏ*��o��lz�m�؅�[��RF�Зe�wx��a9m �RJ)�k~F��K��Z&/L��٥���V��0qOR&'�
�b,��2Ͱ� �^
�hzK��im_�󅨎҉�~@h,w~�I��u��"����"���*t�dy��'�/Aດ�@�G�lJ8F_��È0���焀��3�!N&	�` �V�Q����$�P��x��ArBt�����]��W \�_(f��|2xM���Ng���i=�����4���!(q�$>CF�ǯ��H�̴�>�� �}Ԁ��'V�yNh��2Ë�_�\�y!�������=�4�;�x�J/�2�ᳲ��9�H7'��7��o���ö�~�܈FVP����2�mx��=�����
B4.N��S,z��lKs�w�.�8��2��=䤏h�׳״��Z��ίJb ��/�Ͱ�w�����%~{�-7b�ǘ-K�]����9�X+��m��kroS §$�a��$w{y���-��W]�页J�*mH:X���KchD�P�Z/���lS�N5��7��� ?�r���5pP�:��4j�5k��29�?��3�a��8�	#�hB�?������6k�;N���a����P�s���**�g�G{�HY�IN��gHt��҂9A���<���{�4��a��r�U�oK��"�'[+[�Ԃ������� �C�2j!o�>���8�j`������y�''���7�Oc\%��7�#`����ᄏ�h;[o.�����/�Ryt�}Z�Tԫ�rk-Y=L}��KVJ-�>$gY��!�*\Y:����AiKE��*T���6t�`M�����P���';��?.����\y,�?ڝԤ��1���L��L/9��מ��n	�Ta�-XW�Qq��X�x#���U���R�?���4mP�v�m�?7�P���y��@�WzdM|��g[J4640am�;������y�3���MlWj��D�MbO8qpZ�?�}[�M�a� ݌{Ory���O㮐�¿cЙ4��fDC�:3�+� 7I� Ѐ�G%2�!=e�nMw���g.�(��P�N��������I\�N��2��O­C�H�������]�R�R�����扃ɼ�#�]��L*Y�� U�1>�����6��^�gr�ի,�'��U Mf�17�"��k'��?oױCW94/���D�b��#����'t��&��7SD�Ds���U����k/�mr]WƊ��t��R����C|DL����H|%U�@M_��&:�H?�
�����n4��%�� �\y89E{Y�OB�4P�ؕd��hF-���J&��9s$�z%-�Ft3L�t��a���I�G�T�{��"�\/�t����H���L4<�/�d�{-�&���3��~w�Em��h=�㮠 
>r6�i�������zd���c^��Q�L1)5�q�l�Mk��|h-� ��_��/Y��Qpc�]/�C�jo�%�L
I6�;22�MCķd9��򜴸w��ll{�ga|�hrf�����N,c�rϐƯ��[��Z�A���W��I��IF��!���Xs_�Y�u���x�R���+��n�L��w��O��<�d�K�*w�8Ӂ.�_�����܆�؁cb���AgПT�2�-d���Tr����	}+SA���Ec�"�M�O����m��Pl(h�2'�9ˌ�޶k��ɿ7Jyf:k��e��qn(��a��$1��"�*4�0�<� /�f$]@}S���+��w ,4�������+}cG]-�¡T��:��~^��Ƽ�K�q��;�-2R�F�z{,�Ȼ+�U��Y>ޑ���ȦE���~�����I$����[+h��?�Pq/���)����br��:�*YW���ɽ�����=B�E�&�s�Lu����H�_�J��85m��:���8��U?�Jhr�6U�._Ӽ]��s^1/�2}��E��Y��L*�Y�,���������ޙFP�&'"|j�'��s��X�RA$�K�N�r�۩��d�~�w/y�h�C��?/�T�dv76N��>���ё`|>��%:ǘ������V1��l��)#�]�1DR�o�!h�;��{���p��� ��:����WOmOl�[TPG8�!���䯮�$�7'h<�� ��μ�\K�0�xIy�,{&����d�Bz
�2��4���7�����<K���k�i�������`wJ�W� P�a͡f��.�
x������퍂z�[�۝L�{�q��ڔa
+����M�n��Y�BC�'r U�J�8�p`ƹ�HX&FG����;����g�@�Z�-�|-P?��A#6:���A��iA��N�?��|����Z�fS���2����P�;=�dR��i��k����*�y��i��ŏ9p��w�c�_��X�i��C�{�Y�RMY�PS-�B8�Zh���VX���V�h�gI	ϜA֠��n�[�jw���9�0�z�Q�	�yyw� H�2������] �_>ۣ���50����tNV@�d��5}��g��w��x�<f��?�#s��;�4��ghW�tL/ � ��kl�J�q��IQ�>��<�_�Kl��r�7Z�o��z�e}S�a�H\J�U���,E�O���#c��*�On���M0��)/ڋj���ܼ1(]SH��Rf�j*c����Wyi�J(��Cۋ=P:2���*��{5�5,TQu�T�r������f�ײ��(u�>��.#�1���z!�_��m�&��op���+�<�3�(7]�uo�ܟ���U��:�AŋNK�	�Hsi@�������[t� ��ʵ�18�G��ҁ�\���ƿ��7�DP ~Nᳵ'�}�<7�Py�T���f(��'!�n,�� ��@z���p吵J��e�V�=�U��]Կ��~�����j�D���M��fi�lz�c�-�<�e>x��>E�pg|F����(�/�R٥6�{�<xb0i�E���x�	=-�MVOÚs�r8r��<}h&)��t$����܃,���=����Gk�F6$(�Jr�\�J���_��a���#Y�ON�q9��3r�4Z���=��i�-�-RL/s!��hRkSG�`�7��\G��D��ʄmIӥ��(�$ �9������X�|�SjɌ�87�.x��av�ʿ��|`[ur V�f--Z?��cD!�}w��ǡ�3uK�Küt� �� �����?���S*�8rH�C�JYp�;�b�)
�������d1�;8��G[��Ĥ�*�jqf�@�k���Dҟ��L)�<��"�{�Ձ��in8��1(�b����>���`*_7P�Ϩ�;L��]����mCU��4F�_N�'=F�U#@����s�a�]�d������ څl�Pp:�f�=:���ac;v�Xzzh�O|��s�����a�Jr4��eb�X�������[o�LdA֞�h<�X� Ҧ�l�5%&m'���� ��!�K$�����ZD��3O�V�3��![�a|h���k80�(aéŲB�"D��W�qxdi�]iIv��@�<n@�H���YK�E���q�]�+���:/Ec�i݀
�I�y 	U��$]At�+!�����R�Y��7�؞bA�����$`c!$֩�;��l�_�Q6�R[-9y"l,�v�q	k\ov��OФܵ���Gu��2>����(~L�22tm�#���t���^hF��x�;�-]��?���E_e  H5$0`�É�IH.�ȓ�mD�kf��O�g��(��l��e& �M`WL���x��g�ܺ��o+, �����g�/b,/� (�B��e��Ee�F��^�y��>g����s1
��8�D�<,�Z�{]��v ������J#`�!,�w��Z���;w_C�:���<��Ił0�>K�#E3����gfl�{ U�j)�vM��t��^�W�"��;��_�����hL��#5��RyF�SΧ�L�_�;g�Ƈ~�bnj�-+�<6\mRH�S�}1�'��b��ɛ�a�Uv�E{ؖ~�ؐ_�:����6�8�9�_m�ͽ�ͻ��P�+�[�#��d�����7�����?�^,y���r��%�����_$<�A�w�x���DY�����h|e��\�Gڡf@#�`������ !���<o�XqUn%)��A��G�R�G��,Zqtu����&��[�ҍCx��߆ms����vw�<h�=*e�����<O�SKlU2�ˣ;��9��@M����@Ƅ?�їk#Z�$��~B�~�`�(!�_��[�mrl޴U@<3Pݷ��r-�	�d��8����z�@�%[U]B�مp�w:G�H��|���o  ��>���Sٵ#^�:9/�&��S����<�:�4����KK��W��|ɲ^3�:7���ɍ8F��HMd|e���u��V�o�
cl����(���#�&��D�Ȝ�E#G�ѹ<�x(F��Y��t�VHC�~��)�OmF��{+/��#�(B,��t�>�{��!PZNp�V�d6I_�µ^�����	_} ����:�`Q�ƴ�!B�f�����b��h�v�L�8"�GR��|�:��:(�&	�}����ĿiSq�Q�E�*�R�}Xyf+mybH1�VG�B�n��x,示|�lk[M�Ъ2V�v�N�G�Ec��4�o7�gh3�o�+�	'�Vɰ��j$�1ٷ�����m�\�b\/{D�|�F�����n"�?�I:������	�΂cttj|S?Sx���
ģ�ڤ�Zֳ�39�����a9L�����T'Lؘ��i�z\�N�~��:3�,jp�i�{䓛I4��������L�\�ڭ�]�������z�	��>90	N[:��8cz��l��߫�-����V���7�4&$����+�Tg&(t+�/�SQ�I�E�R&�Ơ��	�li�"�} {5b�a�}�I�z<獄R��0�pzX#��>XːtO'�OE=S�J�]��3������aP��ܸ
T!z9bdfc�=%�ݟ��5��Oi���X{w*cW�r(&yP�(�d{����2�R�I0�dI�C/���4I^75i%,�;��51�r5�5���Uu���y���W[ӫ��	m�K�ļ�B=9�R� b|��;���0�c�S&��J� Ә�W��H��nD�,��DQs���.��$D8H�(TF�6��D��	���@�$r���e�6�����|�r Y%'��.�
-v���Q�2Uz�X���$��̷�U�r4*�E,�������L+�X�<PO@����Jsy��1����>�~9��T��a�q��r� ��\{!�4V[iF?���	p5��W���8/�3D$��pI���� Y�<� 3��Q=
�6�HOUJD��H�j�.@N�k'����V�slYD�n�s��/�}��mXG������s� |���:�D��#k"f�/��[�\RE�Qi H!���l1���骓����9^�O�fj!��s(g��h�gG�(� b�x~�[��
ꋫ��|�~�������o���r/hضy�nn�5vӠD���H��j,,;@*�λ�fZ	PßU�oY�!hH|���J��T���^<�h��i��On���O�7�qv�~���X�$jNꈕ u� H��S�Hj�}kRX�����hIo�T,��@hAOP0u���.��W����!��R�qq�w:u��S��׮�K�v��Ѷl�_=0۰�vp/ J�hJʕ�_����Vx�V�m���e\mo��*�����f�O�҈�L�Ǯ�?&գ�y1�=Jx�z�<����O�'����$6`%��� O���?�dP9K�wi	y �����l��\�#Y�F���k$w�&r����7o�~�48�꓉Њ�\$!��pi�7g�,͗m���%*�t��^���ő����L���������hS\��q	JV��?�'��|�[��W���>�BN��j%wc�>t��t��_	���@��e� �YKB�;��g��`���� ���t�c���y`�م[��GA�a��A�� ���Sr�1�ȠkʝL�Os���O\C�f�x�^���LO��8s�Tgd���򃒱4f�����f����:����\��<��a�(��>�do�|��s��0�+���{�ʉ��'�}x��P,?�n�(jY㮥4aF{����*w#W��e�,p����d��c�Of�z�� SV��[�YP��÷I��]�FP�G�x���xR�����G�B��G�􎚏� #-��<��Y
B��
�W�O�:�P*�U���>m��u�}
�=�0��O9-M�I��Oj���.���z8�I'���j�����D �����.�o��/��B������T��W�g�7W����֧N��;�� �����ȗ�QՂ�����7����]Y���`#���hA��ğO~?T�	�"����0�P�r����`�\�`��!����@��{���dg��,��;6N�{�A�1C�@($�]ٙ�-�.����j
�8�o��	}�p�:�)kO�ɉ�t�]��2��/S#�;Ny '��C���q�w&\-�\�=Ղ�^�]M�:O�-��.9�V"���)%���ƴg6���	x 7�{�G�:��,�<+����>��<�UB�o��1x�f���ؠ����ԏ3Ψ��Cٍ���>�> _&T�q1��ԎY�����8�4.��� #уc�v�u����3zqk����,�%l���[��:kA�Y��%�' ��խ��O
i2�om 77�p��2�I�ϥ����m9ԧJ�s���ߵ�P ne���)����������CK��ߡ4[u�Ú�����#����)r���\�1�a��	���,q�Oѽ�����vV@�a�G/�Q���4U�x�( a�ҹ~>�>0*.x�Z���@�5]�ڑ��F�1n,�d�1k(��J��kڝj�W,��:~i6�RX�|�({��G@z�6�S�O8�BY���i�ي��s�x�&�2�	;���sB����kվ&_��Pt4K|Ƴ}��
�9�x�6�^fl%{ +�K�'�"ш�����QS^�Z�A��L���s��]��ݓ�f���2+H\���?a��F��P�Ըs�u/��z0��v� �]TVl����M��od�d/y�a�װKS���3��������rXژu���h�Ɨ�L��o`��3LM��ⵈVr��A��*6)�B��a_���>�<�t�l͢���4[��x���N��;"]�r�=�b�>%\��>Q���T�d?�v}mU����� ��υ�Cc�z!���㺣fv���(��	$õ�dJ��7o-r�]�ǣ�u%�Q�s�9L�4D��jC[ʳq���|��l�"�����m���� �3$�H|��N��+o&�y��Ԡ�N�^*��}��r�T#������e�7H��v�#n�|ڜT \���əM���a��<7 �m�Xt흃��çX°�ږޟ��������N!߁c�BihY����K�c�NedJ�@~����r�Zd�4��Cx٩G��d�?xhf�Jf,��Gxh��R<�9~Xu!�EPl�8ǏpU6s�ӣ^��c3Y<���r;�uT\�N��4i�]��hKkK)t\��|�ٲ6)	��C_UA5����c̸A�K���a���XQ�n΁����c��Gǔؚe��5��Ɛ)���U��;�*�[�Ju= ����*�x��|JF��`���k#�:�[|՝r���J:Ln_��%�"%	 �t�bk�] W-M�����AπN��������qGl�z�75O1������4��Q<�l_���1x,�]k�Y�����X����t߁�K~~���ο�-mI�b��m�%� �a=`0�9	��VF������^h%B����<�`R	��)c��DM)0)ټ%��G��v��4;�6`����]�����zN��#f����� }�!�x@?��],81�\3s�g]�12��ؖ����âkfr� a"�^�g����o.���k�?�#�Ų~%��b��Y�ў��0��цY�v��Q�}��X���x"^�Q�O����K߉5�ӧYhEM����m��"Ȅd�ã��g ^��K*�g�������ȪC9�!�.�o���������&�r��0�$�G�p��F�(K]���Y���#�A>��y �pw����^ှ�-
0����c5>�^H�n}Х��}�B���A\1��4�#ܤH̔����y瓺&Y\�B7�:���w�i��.~��=�9�U����M�����̦D�=4�H�4��!L�̋�4���2�}���ŉ(��EҺ�ަ��n?4~�Q�~LUw��Y!e�=q��5'CV����O�%�+�l���*(�+�p���j��&a�?4D;��|JwT�Cy
T���	{�+')�� ����Y��J�=�2}:����jI:m]
u��E�
�����3r(G[��B�6S����=���^�`l�G
��,~���4�IHm	��G��W�%0�Y��d��oڎ�g'�t�Z��'W@�k��e"<)��rA+ ������^��V+���<s�����o)2�4��"RP�a2k�D�-5����j mr���!p`�n���?|h��|�D��������t�*�E�Hd�+ϣ�|TXXT����i-�XX
�tMg������H�i����O�<�{ّ��_Cl��{=w�@F7�E`�@D��rU���s(�4^~>���t�Vh��(��w�t�2v��$�h2~�St����:�HX�2��u�g;��%@����@���'>O>2����1"Y����&ZՓW�>G�Z�p���)}�(e���ך��U��#�\��[@�Ah��x�� �+H�
@w*�`�s��QF���Ír�)+	��.�XN��1R�z:"����FY�q���dV���R��іP8=�U�Ӻ���n&#�4f�ɼ/|Svy@��h'c���
�F^f�l��(7Y([�Tקp�Y��ý֦ؗ�H2~;�R���]�މ��X�1��A<��״f!XG>�V���#�{[�
�8_6]�8iZH`�~��0�"�l%g��/�-_�G�ʃ�n'"�`����"$U��+��^�꒣wZۓ��^)OP�P\��}JB���:6���^���B���w��vpTn�dI/C،���ze{A<����;�w�1�m�@LE�}H7�L}�ϖ�t�rTKG�`�+yЫ��T�	�}, �JT�܇�/!�?bm=�%"�ո����cH�a���E�a�t�)پѰsD�-c7��ET��DE��&B�Ҧ����i8O�"�FA����GL՜|{�V�_l��zxjֆ������Dԟ�Ȱ�pJ)W���DM(�x
a�٨��a�[�`��_�Z�bUv5!]#x��b�X�;Տ�V?nsF��4��G~�}w�Z`��0>���%3����q��FN��4;��Atn�G���I��#L_���''2 5��Q��J������:%�1�������(M��	̽U�}��z~_J0�oV~ߗdp��Wk�y�un/�H��5�4����6y����[���|�a9cyCb�B���O���B����ҙ����ѐQ�����Q�9x��+����ڇӬ�{O�z�ӉoMV�(8�V��R<~�gdt|<�lp�E��$��o]���ԺVj-/�A�r�~������0���e+C��ϰi#��w�i���pnٓ4&L��)�I��h"�6G$>��(V8��*R� Kq�|�Y�M�x�)5_�P�|�����k:��N�X�G�!��=.m�̻Z;�+����z�U�=�N?�5�����w�%7��/�r �+�J㫅2�8��($_Y<��P�Y*	�8F�<W'ls�e�y��՟
Z����g |*�_]�aY�3XR�6!5�~�؃鵧@�Ѷc�ER�,�K�d6���2�C	����LcOޮ�E�N%F�e$䔪�F�[�72V�m]Vo��7��o��G��۫��n�X���Ш�F���;�RL��AS�Q�"�=@��l���2���L�KY��]4���yS-6��a�C��J�����*�$�\�Z���)��Ƌ��!]��hmB�d�X�[ټ�$�4�6߲]�~��S0jq�>=d��^�
����~b�`ޥ��4�?��u?!KS���Q��s&�9��/O
@0�ȭk�=�����X����Fw��
ot[v~OA��3H�h���Q��٦I���rN;m'n�?c^�K��ǧ�GC	��;j	P�i�C ?�B��?�7���3\�;o��&Ӗ�8.�T�1����ٸ��P%P�#��ˁ�$�NV�y�PP�?d[*��s9x	��^��f�WmĠcp��@3��\»�5/켻�|`��)e����C\�#&	%�<$ݷ7i<f��&�>Z�MV����>�v�x�^��ģ�+@��WR�qm���#�5u�W��AJ��잠0�$gH�OH�C���1�rL�!{���,��$��[[A���r\>F6^�-'}HC���1�p�%�M��I��3�g��kf��x��
51��H�{MC�D(Օ�◌
�+���q?(�^7�*�O8���Hy��58�Y��Y�\mz:�h��z�&�<@��B?��s6���𴒷w�-K(���Z"K�N\E=6}L��H�5���x���A��ie~F4�gML�R��NpU�:��F$G�D�:��ڴ��ke�!�J��^�E����!��Qw��W"&C�YL���^5�"��g�)�r����Jg�������,9��%߄<�e9���� x��~�D(��0���o<ouTc(�=��%)��j�����y�g@iR�L�4���@����ys���'�1���6?j
�� �h� �~�.�$6w�[n��T�_���7`tU�Л�(�[�4��r8~��!k �'7��:����
���@�#�y���y]v(�0k ���'/�wcZj뉐�K�����|��^��'t\tm��c�[�tr�h��:�˻#�D]]���JoP*=Q�:j^���f�j�;L�3�A�@�������7p����lϊg����f��t��R�'ƨ[q����R�s9g!	�j�6���39������|��Tj�}�*R|y5�h�wC���aK�_��O��Z���"���A��T#��iM�7d�ַ,3/���N���%�T�g�@-�����6h��Y���$�d���.*�7�ovU�B?M#�:&���?�|��	
p@�0r�)S��L��3{�-�˼�`��M�w�~*�����>
6jL';ē�D�y�<��^��	<�4��}M4�~.O% ed�O�0 ��4Vi�3>�Z�Ś���BUi��W��3G�wL����`#7���:��Ӽ�+ 2+�<i�w�=�7ݽ��܌��G����@�6p����Wi^�=���˗_�{�b�F���3y�SX,���l�h��S?�����w�+A�����d7|*��[t�[�mĆ%V�|
+8u����	#��V�������@�DC\���xEL�U��i�'R�O�����������mJ��z�M�v���C.C��:V�djv��>jV����O��ec��O�R���l�$�HЮF��9��Q����˶ҿiT�I�-�*�C�j�#W<� �d9y��"Z
�`\�L� ��I@�L	x���z#��G;��j�j���8�U+������1Z_a����Ң`���N����9��r*�2=�h8����d!�`~g�_2&�"�;�ğ ��� $Z�a�5�&� o�_EM���=�'��p��C�j��;a�U����#v{g������L�=���HV5V���9�bPeu�F����i�X{j;����f4��F)9-Ԁ�7Fl���&���O�뒁C�|�Ғ��i��6Q�����ss��~#Bb��	��Ob|`� �ĉT Vh�/9�*=���H��DK�\5
��\|�C����Ig,�7������b.�+��a�o�C�bۍ��l<��S�B|F���F�㑤|ĢOW��M�F��P�?k�c����ȹ�P������"��l�{�y��qE΂��vm��[�J���52��q� $-4�:�$��r�j𝔖�À�	il� _ @��B���$����EJ��#��ʲ@���S���W������ӹ�k���%y!gg�mXd0�+r���g��L~���5��zj�Խn�۴ֶ	��$�t���Ybv����
�b}a�l� yW5�Ee �3l>���;��E!�ç}�,�a(v�z�:TP �4=�I�VMD ����S�l�L��o��z���w_h��T��x�� W�ڼ�¥c��L������-4Z_��S�!��H�}צۇG���L%��g9�.��%2y���d�����N [�1�R=���j�J0�,�Bt��� T~>����,�;%�o�0�U�{,��4�t��h��f@����tśs ��Z��3���(������|�m�{�R���Ev��ae%��E0`1k 'F x>�2C�vz`T$i��(P���=���	>N�嵜�6O�g�J/�\�F�9� �eE]��o-��,S+�B7�{��������-�%��hS��j��%=o��,�߷��f��*��2������A�O))�W�1e�rU=�?��-�����Gl3y����%��JL�2ȰR�Rn�����0@هg�<lJ;t��������}�]h��I{�3��L9tjeҏ��
�QBV� L=�Sn�؝�C�j�C3�ѹ*�m�p���Yѫ�I�-�zg�gb �"�t��f�)I��&�> ��R���yک	k�1(�v�c���W���0��^g��Gl��D�1�L$����f�ͥ\3?�o���U��b�Y��	4�P�94D�/���
���:;�*��GP&��Z����S�|^@:�>c��Ĝ"p�V�-��,�(G�;�D�;/T�u�yJ+�Z=CF��܎�?��X��2��d?���[�e��?=5�_����X77�լ~��D���@ W�Fx�^��Fc8/��C�r�����|'$�?X�M��;& �s��7�۵�l�z�z�����r�0��@���R�5A07���D�7�&�7yc�C@�;��i�/6`&4�����BԳ-������G�E�g�)/����#J{��~��҉&IN�pY�A���|�-YAB�7��UNvb�TS����#�]K8�kI~����2�w�Ev2b�QQ��zsYƇOi"ϵY�
�̅�ó��'y� �
 z���;��lL.��+ۣ�B�Zj0�����KV�@5:��PI5� ��+A�}��̫,V&�!v�����-.�@p-�޺��]���F���=:%w��-%�_1����@�;8Z/�=$���+.������b�3���d�tǩv���0�_�,��|:]�� ���ѲᕾQj�6\�nꢁ!eV��V	�^#l��>�F8N�,��-����¯D�^1�j��6Ø2�>w���DV��nO�=#R;�����d��Kh�l��^.���+z�3���9i#�����Q.���%I`0ȿ�>���Pǝ�
6���.#�Y"K�+����u,ˋec�N�����m��b�RѤ}^;m>ԇ���0�
{��f��������8�B ��;���lk<ʑ;�����脞�7Uj,�Õ�aj�)�1Զ4��[nm9-α���~g��IJ�'��� �S/W�pn�3��KcC��I��r�<�=���^��|E�"6��a����o��ݺƜ���BMs��z
&����ux�I�Z���&�氬k�G"��P��������(1P�n$�?ęc�h �y��@𯩚ق��%?�ς���N�8��YP����!��]�`�U�
��Dc{P�P�X�-T���Rv�i�$ZWm�=~���W��}�V�P�$P�'Eg�>���e��ej�C�����M��!���q`N�64�o_Oc�s/s�v�5�����2���g��|���������ڴ���N�y� ��o�]�,&I�q��Ӹs(]���n��&���x��"3B{�ԆT�]��	x�!��ղ13>���G{O2��h���bU|���= �
%������ր'4���I�7���D'	�IKY���}ʛ�����fѵ	��>�$jĻ�����p�B "�^�F����2��1�˿>tns.!2�G��
b��qn=`�)���Ǥ�q��hn� y ��7��k�{6D1�@$7D�`(�?D�8��M�h80�cz�����ō5�m����mD�*j��!��K�rFg���n��T�D�\�w�/=�W53@&o�ec5��u�������C���4P<+09��̚�Xr2��*c��?&���4��E�g�b����5|}e��`��ط�ћ��F��b�H��L9�?:QpM�3Fӄ�|G_mԊc��&YbbX�Mh���ҵa}Q����cr�a2�H�`Ğ�0j@�Z$I��ƁT�c@���qf�3�G2��NTj���P�`F)3匯p�,$�ñs\������:[6��-I�����.C�
ր��N=f��FVp�j޼;"�̱�ߙ'>v��T]�v`��47g�0.,m9�w[F)D���S�N  �*�@��WU)��8m���#��C��X�.0�w
����)�$����,����>�5�E3)wD����g�������)��������1��YH����P%����xB>k���h�����3��)!�u��9K��Zɏh�٢JM���B���ʎ*�3d��(gr}�0��< �q�¹z)�}�b������W[�1�5���iɚ$nWFw��_�"����:�����U6��n������j�/�!���̆�l��!�ɺ���Ty��7��E���\��q��o�
�P���z� ��A@x/כ{?�ou����m�C.��x�Ê�}��PB�E���!�wp�J%��K�u.�����>|z"�� ���,�-h��>҅�׍���k��:�����a\���'˰Ɣ��^�A��3�EѤu>��;^;BSH���pi~�*�V��|�3�c����p�
b:�ݯ�/'4<��D�7o��~u�%M�_���(�Z��u�p&v��N˙R�싿/A�3�2��dg���+�3A�}�c�u���z�ZQi�ʌw��U�V]���6]E�щ:T�TmQ!Gb#��	�yyl�����9�#�b�]&:|��������1���sQ�'��L�fz<{��%w}�����ҷ�LZs�V�}�7�7&{�M#�,mz䳶,]c�].+�*�U�z�p���9ɜ�^g��"�MJ��Z8�J�:F+�<�XƖ�D켘�~3O#�Mt��z���3dG���KS�¼�������}<��d��H����bI�i<��'
��W��"���T�y�ђ�6�B!��T�V�����Yɕ�\�h-p7duS�^���|P���������`���z�!������Q�|��r�k� 'Q��7$�S�[��(U���H�
&�Ւ�o�47�kck{˔�S� �48��a�g"2s���:6P�`$����8�۪�l}�h��D��u��}�F���"���-��N����6��  M��-ַ~�A�����U<���U�������X����#�Qh����~�|L���p��/V�t�c�xǪ2>@*C!=�	���N�0߄4^	S�T��\�@\��M#e�����-�닌����k�z��ܝ3yA�f��$
M�6	�u4�[9ݹY[���ܴ
/\z\|��4�H��A)\�*R|�JS5�qW�#^9��<(j"r03X����*��4�NK7]����r���yz�ɸ,�Ղ�6祵n� �*�F�kO(���Vr�@*�e{�f�y�6f�O�7otn�dC�� (�%U ٦��'�� �Ij�s CH�jCف�-���hַ�{��+a�e�	����T��]T��hi�)8�y&t����6�9��|���M7-�ojl� ���4�t�S҈�ܖG�D+��̙I�D� �kTFM��Oq��m;|�������p�Z���*�|+� @�wj����Le�"j�~��~����"(�����S�fsZÊsk0n@�٬Y;7�X�d��2g:�k�X1$|*Â"ק#��i�u_�T�q�(���4�gM�|4����"�硖���]�Q�i�'����P��#�ќ���
S�c�1�z���]��]62D&I�z����Cҍ��Y��(3����н�LxԹu�5A�%�*1������wn�r�uX2�,;���3>=v�s򙥵
��8���POjz�}�����~ih���S+h��wޢ/a�H��ǡA�|�?r��X�Nq21D�5����ƶ���)"�H�{~�g���@�+�L��u;>��.��g�^?M[�j�%+��Jo�_��B:��7Xc�*V O.D�h�JgS���e��b�|M e(K��:xi*kyr����RU���)�p�po�i��*J����t �Eƪˇ�����!2Uc�ʒ���FxNd+<N���	2s
`�a���)��z���^�'�;D����ً���3��`d���<mfq�t֑&whp>��=
z��Vy�e��<�;F8~nN�t+�id�k��%�Ol"����� ��0�߽ȩ�-P�+�n�uf�ZŞNɶX��`X��%�2ϔ�ly��po���nf_��b���	������H,��,1�v(�ax�Gt�T��ϴ=+�@(@PCW�Y�V|0�#s ���O��w�W�:�D�GW'�L������p��
Z��U�7�e��޲�uA�}	y�»�{�~+�L�`iL�"�	��Gt�.J��F��L]v����nWs��j���@̗B���*:q�*�s<�U�l�*��~�:`����R2~�)�xק����>M �D�z�[Sι���F�מ�_m�Ȁ�sg}_F{�A!;�X^Y���B��ZH��be��Ԭ�씷u��8�Ѓ�N�fla��y�$;,W�ŝV�x�G�4)6s��w�O����y9Sf���{I'd\����d>��������ؐ���,ĚQp��ʳBI�L|祧=� 8�齺����� ���1�P�/c�o5#{�s����=|�هsw<-��Eܽ�Y�ژF1_L3Z?m?PyN]o6�	�Haݎ��S�+ṝ�������~(H�&��Gо��b��rBӾv �йy������A�VK��?8[�i�N�a���ٮA��z
`�SO-�mTDQ(��P�&$��j^k$���<0a���r�h���]�m��A�Oc�:Q����<��2�x�. ؈��A�u^VWB�fB�1gF������?�K����Ga�^ʷcz�N� �P�׏�t�qr��߷8���V����y�m�`�ۿ:9ه���?DL'8,��o��l~�b]]Pz�.J{���8�y�A�Q�#[#s��C�\o��+�^+�w$=���c��X��/�ǚ�VhEU�Z�u�$�\�U���ݞ�W��3�������טRBj�>�G���S�F.�(�ed �����K��^}-���[q�HpˣG��=�d�Vp���l��$)L���FB>*1����l;�'��Q��Q*�����LJ$��pMS�g*���q�¼��\	�����=x?
J�7����y�ga%LF��Th��SLb���nxT�B��:!ԟ��E�b�W�+Cs�zx�w�8�:tu%��:$0��B���ʿ��w�o�!o����˻0��@��>k���>�M���j� q�b�O	P�t����l��m�̸͗��ܮ$�{k�$����&���{�T���b��˻de�[�0��e����o�W�z���kQ�ɦ9f�MSs�y�ԟ�j	���7VĄ�!�C��0}�QG�A��	Z�"���!�m�
�(��?�����+��M��s�R��%C��{jIIU)���6]���[K���_�s޴(�$%�H\�P�@�]�8R	ĈW�ˍӨ���>��� u6�ުJ�a����q��FԔvy��y��=��X�Q'�-?B���sh�Q�d��Uj�-��J��w���Z��!��S�kv�oG�,Jpja��+.�Mx�㈯}��7��Opǌtuw�t珋��8:�p�Z��l4�j��+?){�槶�7h܉�°���gY�v�9]Ew�����شa�H(���Y���)�'<�C]	�H��l�N�0�q}~)wPE��{����#_ ���y�5�+ �N��cQ�QC���
V��L��Ӷ�^�^�Y3�?�Z��#���+�*�G�k͏�16^vWMw�a�~��R���MT�d|;  ����[1F9�R���c�����3�&�^!-x�ElNhM��C&>�Tb�t6o-$����WR�y�5�^�n3`vC\e$�vp��h*˺����/�����G�U�?>Zo�O4���J4�xI�&^��~��cy1�O��������3����8�j��e���L�W/{�K4�#k��i�R?Q��@�]����(�8/�d1m78$-=�ZC���s���*6��@�a<�N�})�8�[^�ؼ��c�����nD@�nl����Rk���˱�P8-��/K�؈]>���s��XB���0�wU�̒���gy��߹��J#^���U�6�!�j��``KÑ�5l��4����
7�,/*�F�%�9�^�^�U��"J�� ���_lq$��������&ž��˳�Wd!=8���y�[� ^Ѽ�����\�`C�f��^Q���#3���w�r��L�0x���a{��@���p5�kf��E�d87}�5p�0���J��Y�66N���I�����Oq�I�T�`@4���
$�½�o�!��/����_�y����z+��G��ۆEF_�u��i�bY�.�=f45�r�F ��R}��H��r�`�q������r�:�'O���1�)��Gŉ
�=M��aW�Կ�I�@�i�;ϙf	` \j������	ӧ��E�(�Ih���#��ȥ�I�/Yϣ�X���f����<0'��D�����϶*�������~���(:[L���!<[r�x<���ۤ:-F����s��G���uc~a4F2I`�f�ּ�br6	si���ǨY'��0�3i�g�)���㳌�����|���̋/�l���}�ʆ����Sv>�7ͼ*�(I���������K�v ~�,6���%ܓ�U
���[�픗]�I��=�Z�5��ŠS�:u�bmȳӣ
p�p�D1�߾�{J����p������݌[��܁*#�}�\f<������.�3����ù����Pą�
��Gܚ|/<[D&�+L��������Vk\c�����<I3�s����1
�u����v�d���nD넼�42�>�Zq$��)�QΛ�����i!L9��/��[����ݻt3��9}�C�P�zN�Y�j2,���<5kS����/+=�-wF;l�������@*{�j�~�/��&�j���a��3����C��e씐S���xi�&�A����հ���6����I6=!'�omt�?n2$���@G��(t���t�p*��>���K���'.���M(_��� �-��9�i�*�+ٕw"t|�k�ͱ�CM`z�N;0��n�Mi��E�j�L1*�)����5+��K_ %N��:�Ψ���JnuL�/ұ���f���DC�ytu��\���=+�v�K"菘o���������T 	��h؉O�Ei/�9���^���ĭp �-EWVa��cL�p$�>�S�Rd������[�������!��� �~qJ΀/Av���1�^J�kZ����;r�$r��GP�D!�y?�ی����{\Vy2��ܸv�w��]��}\���&%�|������<�I����B��vY�-�\��������e���n[6=H0�8���W��F�*P�^db�vǚK�q�H���m� �1�勇�ar������PR�䮀�0��Y&�+WlW8�!����@���d5(ޢ�W�V��(M"Tvm�1���IJc$=^No�>�aKܫ�,o����p�-%�#�������c0�JƷ����Ƴ>�-�j��_mǶ@E잇�^P䤄v[z��������o$��sl�!�ÁF�&�V.ǳ���A�3��9���Z�n!B�c��i0�Q�0��gsgk��Z�)r�[c��V,����i�Ve��Z�Na/��/�+ĨQ6Gʍ�0��E��.��Mޥ$�wB{+�Q�O�JG�PI�Tc��n�Hp��ӕ!�Tr�����
z�K�L�6��iC��=6��i��{�la�s&�>B�G��/����/a=ƦHSͨ;����/�D�o{W�O���V�7���ӤS��y��j�Z!�^���}A� 8 @Q� #��ǡ�s��װ�tR1Z�����z�!f��
�E���Ю���O�k������e�A�����+�]�i��fgc<�J��X[�����qo�G�F*�0����X5�{ß����@�\q�"�E� p��R���v�U���p��u�\���2�������݄���p��j�[�t_X/�Rb�NS�ɜ ��Yy`�}��*_�e)�i�$��{}�~�1#���n�f��ɗ×��<��+u�-!�<&�,r��`x�@�6����.�9K���%7a]D�zr$����9������AyyM����ld�d#�y�ٔ�(AC�"ު�i�N��:f9om�W��xY<o]�͙�+\������؍*���S��.��'}t�~R%i����ފ�U����gw���d1�s�9��a�#N`�M�0��Z�q4�3p�r���L��p;W�g�o%t�uM?�Sk~>�%�1�O2��g_?c�C�N�D�=�	�Jp"������i̛��I;�U�E݊�Cu�$9��0�QA��M����8���d��^i��wuH�ΰֺ�pO�H�β�,N��x,�COڮ�"ƃ���6����+`�f��V��Az�$�x(jW_�U|�RX*�$���Rk$��}Ĳ���+m�Yp��{Gb�5냓�1�\������.�����+<�TT?�L�nezs��}�X�')�9���;�[�����2z��^����E�Ī�U�^���q����T�MVI�lW��W����ye���T�o�,Tu�W����N��nTh�B.��3�N�<�
QzCf_���T^ϟ��B�V�D�!1���Ǖ,���Z�m@��DA��;g�rP��$g�+>b_�I?��]c����{��uw�G�>=�L\A�����qF��P!������cj%#/]!��q魛���U�&pK���u�[�X�d����f˶��y���M��1�Qq�/vj�����cS��C�E�D�%>��6Lϰ��I�M����?x��V|�x
;����Pj�O� �U:I\�>ʆO�Ps�1�p�2�cP��Ka�ur?��P�-ǽ/�=����z�n�O۠��G��>B'v����C���n �'[�c��A��2�(�)0����-?EP���S7E���E.�؛n�v3�ؘM�JT��&�o�_GFV���a'�%ή3}�N��vyl��<�O�6�K�Ԕ��M��~��B�Zz���n�8%�e{ϊ�~�^:��Ҵ^�C��"۴�D6�8<B��5�$=��y�/p�;s籃�lSn! ]���;/ZZ�*)�\Y�ù�~Jq��{��ա��b�g�ٮ݄^h4�큲�=���50��-��'SV��Y��U�'+3Gw��79���L!�pC2�P��R����ʕ#)�MA;-M�l��l��Y��|��@z��.b>�c1��^���ē54]N���c=��ٜ�|����/ʼ��֊�vJ��d˶�~v�%.yA�w��tV��E���jz÷^���mP�T�[)C�˵����[���eV-���@�������eܐ�k�z �S1bÌC��Y��z�O����F��ub��dd�!�q��>	k�wݔ�s�b~��� ��	f.�C'�Ι�:j���r�����짉u��^��m�U?uO��^�����"��lE��?߫�~)l9��`}�'޿0�����ޣnV�f�<���Z��<�˷�G*C��df}*CO�z��j�ؤ$VZD)�cha~��Q������t��!�������_{�̧��P�^�	>��#C~�yO����4�ɃB��~���;�[T|Os�ʉܭ� /�%~��7��h#s2um�w�����EɄ�|�z�"��1	�*�I��{���^���(��GA��F4 q�uφ���F�7�K�^��^�%����Q�PȞ�kr�J�>�Cͯ�� K�
��.��)��Z����W˼5Dn�F�����,���:f��f##l����4�lx�����b��TYV��v�[ٖ-i�
�i��`��f�����1/�dӫvs*H��?��:VJ�Z��WΨ�6�"&�Ҽ�*a#4��	�qMㆺ�L�#�x&!����ah��S�ߢ��j��k��dõ��]:R+`�hv�����4 ,���@0V�>B����-^W��{Ob��_.ii5l�b��R���SjK��H7?���vCݬ���g��L9!^0H���=�t[�+e���.�U$��į�&�o!V�*��)�%X͞����I����?�b�l���F����uN��WSZ7Ϛ���?j��w���#���b�
�!4
i�Ĥ�q_]�E��������7m���q˶���93Y��+�7�.�JxsfD5�֢�u.�L�Y&˛��ר�_������v�V󶇱ۻBbO�%	�p/b�8��W��(dmk�2Sl���aw��Ӄr����%3��C�s�`4�Kb�<ք�������x���o��x����)i��C�JI��|Z0T,h}�c�S{2GW˒�-�s#5��e�i-a�J
�N��8�~*Pa��x;�m���A�N��Z�oɯ-
�@�KpQ	�3����cbP�mv���p9=�{b��ɽ�J���\ʣ�����K�[��h`�չn_UC�j�.}h��Aߥ/Ƽw!��4r��b��<�ˑ٢sD��I��#mZש�sR���ɔy.�����V�Y��Y��7[�:�^-�Aq,�ږn��%wȽ��,������W�Lp�\�.�o؟�^0���I��"$
(���5�>�
��D��\74�:2�2�����wT��Q�'�9 ?�#���ӭ>��F�8�$f���Ѐ[8�o� ��ӒTx2'A�-�էN@x��]����lO��8�A_3�M)�z�W�L�<���\�s�՘@SS��wΪ�̩p����]��b���w���̖A"~��Z����_�o1	_"8�T���ґ��bL㞲xIb�3*�ʪ�0��D1�ש�7��*���*�F��?(_?�~�����Co`̿�"��}��kZ�*w"خ����:+�3pv���ގ�i�Ú��	�9-�j'�}ʵG���w�θ�+�M�^ѭ:n�^S�j���X������-u'��l1�b$D�.��RK��X_���Su�T	#��N�0E�axj7��:|h��'���SX���z
J�Q��M�f%�5Z913F'
<�U�8��Ǧ}����N�>$v�bQ��o�j�+�J�Ƃ�,��P�_�+ᖩ�q������G$ �8�r�?�;�9�)�~��9d��«���V��ḩ�ߎn\���|K�:�i��ʶ�g��s^m�8du{�&<Æ�	9�!z�!3�1�L .�[��6��!����09߅���
�+,n[�����R�\@8�L0o4o&m:<�
2h�+����RJ�:Ktr_C ݧ��ø����5Gk��~��I�L�O&��-Q&��2_}n��Cܧ>�6�en��bS�=�h2)�<�n��:�?�S�� ���ؒ6ef��p�0\5�~/���y�� ��B�.D�<E�̠G���K��ؼ���U�3��)��S;g ���q��L�� �^�|��z��N��`��M���[�GX��lhI4(C�۫�b�Fs	�(�M`s@���G�~������q,��g^kx>���CRUb�{�[��9�l���dF})%Cf��x��|�bV[��?�����:HF�=�F;�̣�[q���kG��/�nF'�VMR�i��0W�S��o��?�i�v�sk����lu ��J�aG�׍����i�*Sd�t_��nwSUbq���PX�%V�s��Ռf|`�Z�:��S�w�����ZX���=��%�q�/K�
��N,���jzd��=��LBN ��Q���G�~( �Uȩ�p)KH�Vj�M����!�\}��e~��s�uB���N$6 h�&˳LI{��QtP�T���l���{��bMS��PH�+���/���-�j�,��jP�8E���p�o��i:�}��l�$��Qe+���xF�"V�[�!UM�n�+�CtʄԮ'���r�n,�����T*���GiZ��3�����=0<��%��k�}1�>���!�2��i�ucuh���;/&�k�'wz�^���zEEA/�Z�D�䳭���.��^>�=��~FB���6�@���K�����T*;��fXg�鷪+�d�F���x/�o���+��Z+����=-c"Ă�9��-lE�kM3�&�����V"V��w�|�r��sg,�����į�����HW-����e�J�t����_ȩ ۀd�0�hU
��=N���<B��+t�~̇��j�ƹ�]�8�S�.�u[�Js�<(
�!�Y� %����DB�����s�SO>=��\@{�Ѯ6EnM�~��V� 	�-��KGS����������t�T*bc��_9jڦ�gZ�u�h��͔��mx�n��Yh9�&4?��e�Ɏ��Z�����i��A4g+��L0�C���*ؓ#.�F{{�WQ�nhmcٖ�rF��/��E]�3��_�����x��2��9WU2�GU�NҤr�iG��T�YM�L�ʈ���-g�P)���3��J�TS���8�X2jhvY6=��mSo���Z#JX��VQ����-�q�*iN�Ꭴ�&�p]C������&'G�jA�8=jJ-Â�&,Ĕ7U5~�an�W�jLB�=1�s8�bc/�R^�8լ_�����R�'�U:��Mִ=�2�GG!�y1j�~-s�>œ9<���-oi���h�{4�SLq�k��hu�V�\Q��PNk�s6�ɶ�Y������+6��/���Ӳ�'`oh��ea��?�1���w�݆{8�qs#��Eh 1^��	�nA�[�	�<�[�5Μ��ao(���eW��T�R��1�svl���HNz| ���//��޶۬k��b! x����.�Ͱ ��ཥ]�^��_׼�<1�]7gc���#�3@��tL�b�~��OR�Rֽ�˗�������}ͺ#k`�ŅNHkSb?��1!�����IkR|��"��dR\�p��KS��q�y"�2��xj5vXH��4�7���pk7\���Wk9�u*�uzȗ��3���%lDȦ�p���f|��αUc��9�U�7�%gbt%����[��6W�E���� �a7u�&�7�s$>#9:�nns�Њ�
��(Ijz��	`�9�ڜs�W��j�B�����=^�+�&���p�O3h=",9�
�z���#����ؐц��S8��pG\2M��k���@�^�G��"=�zG�v�&`��`�+3_QB�E�0�.|F��s��FX����s�K)K�e`�_Ԩ?����$(7i�
�c3�%�1vF�
�<ZL��E��3�+��v���a\o7O"h��Zd]4����\���_c�&�+2�vX
�n]�dȡ
n�3�{�[H�p��!���r�( ў�/�S�e���d��4A��P��^���$��vh �w�Y�0�"�NS���z+�� ����r������[�r!ke<�!��kƌr_X���q�2��1c4�Z�d�����m �`
)��Mף�MG�E�*��j�;Y�1u�B�����k���{�������� �B�5td=�h��T�a}�T��u���͋?�cpEղN*9C^=ws^i.�6�s�>NDJ�Z>IV�e=
��н-I�m{]\�$i.��Aj��ތUK�p���DKJVb�/��
��c�Qʪ8��N�f��>��� Q��HO~Ӭ���=����g�EjU��S}����!�A��1�����VA	��ܲ���H�mF�l�.$����:��\r��g����U%�I����*�7 !��QS��{}J�a������m��u4͝���d����/pD����L��O�*�X�1�|� �%���<��m���Y���)/M����*�T�`r�]���4/5�PXf��:����}6fz���E�M.[�E��]p�ۀ�!�.4Io�X���w�NP��*R�\B��\T�=|7���%r��v�[�ռ�f�4
�J2��zM7�R�|�>����a�8��߆b�p��x1������J�)��yͩ�
h�pn����K�S�$�I�lmM��nsc����~��� i�p����_w
M���!-27Ϣ#"�%�|���I	Tk٢�G�1�3a���cTUdt�_�m�+=s�� �.�:T��?�㬥.u�7��R�ƒ�����Y��^��BfE�=�^�K>�� ��[��0:薓v}U�Tj8UuK� ͠���l�8�(]"B6)1�����ۇwV�)0�`���5E��E4���u������oE��W�Ͱ|	��ڌ��dMe|Ш���1M}x� Iz�h�a;�Ek�E���mD^��t��h3�����>F|,+�^���쵳{�}�쿱�<��>��a)Aj�s����i��yX)��qm���8�|��QQA��^&A��1w�I�3L7�Ļ�0�|���X�jn�^��F��+�
J�[��XG,��a:���=lO2B"!��>d�����w��50��	D���^9c�naǗ�$�^���w�`�؏
a�_�ةA�^�yb9h��UL1B����5�?sw�*yZz����?�	M��i�7�����Ֆɽw��A�.!���E~��}(*`f2����)���Ĳ���Dx��b��]��+W�8Yhp�@g����ȀWD�X��L�MK����Tcb��!/���>K*(�Ɵ����H��-p�t��gɑ�P��rp<�z�ʦ�^�&���1v9��L� �F��J��s"˗9!h�c�"n�xʊ
*0�:����N^�b���z憉\�8�T�r�A��j_SK��U��^2�	��4g�Rxy�C����2�	MI�dJ�=9���|L����qi�y8MyNq?�WP�h�ǚ�U���,tgx���B�L-���ϹF�Qpܔ
��>�4��`�\^ P*`D�������dJVĪڏ��T_m�dreb8j,�]�B�|��Ӣ��c�80�n�X�Fm���$-Pv���p⭇�f$��v�{2�%yT�Y�Vv �1�Xv:YЀ���31G&�u����u��W�ttad�%Ԓ���$�1x����)�`�hҋ �c��/�H햄
�=���k6�����Ѿf��>�ˑ%��*�M�Λ�q@@%}~�;�B��#Gb�pв��o�L5Aw���W��b�<�%N{"wO}x��!�yq�hů�S�0Î���~�3���yU(v�L��#�yZ65�CG}��h�)c� 8{�<���p��Y��%U�hگJ�-���WM��dA���a�z���,���pC�I�#�p��|pt�	�����9����LS�֮ 7E�,�������L�Jsx��,&?YXF��#�OE�[�4Իա�O6� +��-Gp� ��M���	��+���%��+�a1#[��EV=?{�+�pTE�;�<�.�$zd����Fߞ-=�;���1�u�5�� ���@��\��/�Nܸ�ʄ\&ͣ�!i�m���7ZQ��Y���/��|J��%G�7��y��I��p�WJb�4&4��腁c�|�Ũ�rQy�C��:��>z��,����ڐ#�٘��|⸴��&@��@b�m�TN���C}7�Յd�G�z��g=Ҏ�5�ȞnZG�	�hƒ��w&��YdJb�1��S0p|�VR�qB�:�MX+	�j���ґny��^ՙ���we��=ٖ���+��#���ǫ�bQ�7V!��;�_�ƅ���.-��ZDB�bML7��+A����ȔL|�;�(4����qh�UH��$�;��J���f��mX�A[y&�a�q��4���g�g��j�8�2�xۦ_���K���n+�#v�<�Py����f�I��B��V�z��Y�(�$vn�[N#����l�A9�E�r��|�tG�U1D�4�!�/��.S�f�����7�$Wp򥺡�{�^�z5����{'v�ydw���YA���ʔ��~����刡H!&TU^��j�! ����z�`.��-�o�(�!@(��볙뙊�2��t���.^H��`
gױ_�~����ָD�UQ��\��>c�#�����Ad�vX�����N�gm�ƌ�Hfh���������8rnN_<ڗ����>/�!��D���le�n��3/�ib�����5�#�9��,��s�T��@�%1.��Y�tyyn�
�>�	��h�]QHktiz�/���Il���0�֤ʆ)5ivj�)gS I�p��!�*a��ߤC�Ю�ڕ�LŻ�� �����H E�`����w$6�'6ϡ��'��Kqj;33���U�> �(x��㠾�D�JU��U+ii��<�����L��c�TW��!_@�i�5Z.�R0#�X����S�u�r�	Mn���A�eK|�V�dNx˶ؔ��������iV�����W�4�duo��ÚRr_����U!@ ���i�$�����q�[�:[$lom����Br���3~P��k6�CNn>�D���PW�]��5j�z.y���pA)�	��N�N�A�I�HS��<�XZTw� �� ��Mp�x�\_�B�/��-�Ky�����ې������m�A-���C�N�޲&����¢���'1�0�$���3��8�]3���m �g��Z�+y�pE��P���e!d�e�^҄�6���4d��"�l�	�L��j��9�B��s���6�$����j���<�����sp�m�z?]� `p���0`<���;���S��]���v��e�ZViDs^��?U\9Ȋ�������ӛq�ZѶ�;�SQ�M<�+ٔ��
[cC�:�:�4�y�Jl{�1�3<Ox~�Ж�֬���Q9�Tvٴ�*�r��φFʳT��\��f�����F �Ql��jND����T�~��w�'�%���h�,T�F���"%�ԝ���.~ԧ��Y@���oJ!y
7�.�&�L�^EmC��@��I z��ȭX����`���}�;h\�^�r������y�8��ē�Z��&���x����>�	����rrs�S@��t0����-�a<򢒳 ~1bȏ����|I XR	<d�c�b��s� �a�Ѫ1�;��.���d	�޶.����x�H�}�9ZeVJ�g�d�Ǎ�	���Ǉ_��C��_�z'<�b�5P��i��־���\+eB��z:޵{�8x�{���ZϋS����ᨒ�q�Z5����E]	�������1D<�:}�83�qý�Z?I^I<'�� ��x~L�s3����K�n;N��P� ��:|�k�"m�s�-1D��&X9u���0��/=kg�Oӷ�u"�>H,e�u����-9�u��_j��|"��S���>��\��^@�����B��ϸ�s�1?�_�>���r�q�<��+.}����zV���al��/F�4�.�qŻ�	w�U����Z�#�J�i�}��Π��N�s~0%<����[�!�X�R�[���L��9We�<�<X���F�='����{�¬�$��7��������))�� �=�8sFoFSf,Z}b��h,�;��J@�],�q��uR�[��N�f}�nm�ttrg
�-Uڊ@>�k��,����z�&/��;��i2�Hx�������0�+�} PЩ~߻�i��k���k��(�C>�l��8��x!�-�bw�tAX�zE�q<T[�ӌ�\�0�W�'��׋���ue������'u_�0OR}��j�hѱҲk�	���
T�Iu}�x��ɱ�<z�Rt~
�[�����6��`�]�L�^���T�}R�J]�칗x�@g�(����_%f��>�j�u�PmU�E���b<�����̞_b:n4C� MM��r!
�� �l$a��b&���B`	+&J�_u³ƿ�3x���>u�����^Ž<��I ��k{UK�Qp2)���u��֔�a��1����;m�,��	!ɻe�`�1�Q�'xK)#^��[!������L&�rX�u�F��1�Z�����o|���,UD<���Uk��\���n0;�=�����/gh@~�����WdCY*Y������0g�I<����h����C
8����%(G��l�;n&{y��z�䞼{�z؅G�,�k�Y��o��7�{G�|�&V+Cr{�,rt�.l�D���wQ@-�u`����8�n��[@��{n��o�'j�W��t>͕>o�Ђ_����A���@S�ѻ����<�Q��N��b �T�%i$�Ua,�*�����l�wX5��p媕�|<n8�;fe�5�����t�����R�����t+T�����6^|ݷ �����5fV��þc4��W֭FK������W.���6��D�G��hDY!�46�2���B��F�����4JdI%��Twn��Y49#a}`7���*Ž+�:�s��Z7��;�s{GиQ�2�m�Qކ��p�m��3�x��2O�T���V֫ۤ
s�������k�ӭ�=5_{}��1]�>h/j0?j���͂2]	w�$g����P�R�����zܵ���J/v+(n8E4ݶ=?z#��R��i��� �8�ua���X�Z���bz�c�<Uͪ6�m��0D����a!r�"���Ơ��}�\�7{k(g�;+Ѳ�k���uCr��wDk�|�$q7�ԣ����آ��F��۸��g|r<��V�I�Ѝ$�0��{��ę�+�6O�R8�Q�^L�b�W���`o����P4�{�I�([����C���A%����Ͼbz��Z	8��,�ptE����&�
������ι�e����^�Ы���uO�K2�-�Y�[뿕��83���'�Dٞ��MT�����a���k�sѩ2x���t��Xw�V����R�� �tG��@(�$q�	�O�����S�5]9�m�'@Ý�ˮ��*/�GMӲ�t��_ؐHc!U�RR#O�3*11/Y6b�ab?�Sy%�kZ�-	�#�C�w�'�n���������o�9Fs^�a��]��~5���������䶥	�o�w�-0I��,o�"28�4�[u���ont&�8*�`)�}H�VS3e��`5r�6}T��ڶ�x�{c�����J�Q�[�Q� ^_��r�^����ƶl����|�
�L�w+5%�5	�����2�[yw��c(�+ReCA�o���)4P�4�s���5��F��i5�J ���G��8.����B��Rg�˺���ɨ!�F�ԏ�%B?>ڇK���`��q`��n�}�\�]�2�w�E��-~	O�  C[��|&���X'!P��QyϹ=�r%�$��ܞ�o{�'�ۈ���z�
�^=�$f��b�	b)�������KSkPՈ�����j�%�.��ǻ��2��LPj?����l?�-���My6�)���B�mt��!�� ǶrF����f@H�l!�ĢX,xK8������l|�l�|�H���Z����c�w�(;��yzذ�e�w��s�M�!<S�]"�V�V��3f�6?�uޢ}�ٝ�A�Z݉���!-s4d��f�f#Y��&�U�G%������cȹ����#����#X�`����C��W`�u�
s���^�#Ѵ~�]��m�ۣ]��	��T!5��;!���!��%aե,ѳ�+����HC�c��n�$�^�Y����y0 N蔿�Ä#G>q1����K�x��\��V���Q��<����6<-l�	�D?�z��簭.���vqP೉�	
w���nŗ����5MXf>(;n:�Wj����9�"�ɐ��X�h#X��/t���U@�v;�J�+�	ۖ�ɺz�%>���� ��G���ib�_��w�/�\<����/<;G���W�\?��p�
v#6���BosD���p����)���w�����j�!��Ѧ�)V�A&f^g
��y.����fȹ^�ؽ8	���	��c?P�sC���}�d��+�>)\9�y:���\�	�@��̢��q7�U!Ĉ��[��u�V
J{�ه��$�K{�;
�&����f?�o�*A�ߛ�&��MD��cǇ+��nsE��pY���u`�UiM�f5��}��81ߤ?�*� ��ƅ�����م��⫿yK���#����~Oj{\cU�8�{�(\.,�B��	�5C�֖
g�� �ʔ����R>=]�Y�uز��.��ԕ&���;��o�~��t}�/CIߴUJ��O��x�m��=��w1��*����
V��"�B��X�畊����q��r���̸���L\ث��>��  �sq��.�9�<���e$�i�q�7\�r�p���[�?��g�7~�P�~G4��os�l^���HuSq���/��xO	��x)����U��ɾ6�ʾ*���L��~��6.��`�m���!��r:``�t����l/|��$�n�p4�e@��N�Aj'�/.8�=�YHP��3���z��^0Yk[�5@W w���:y�%7���H~�v�kM�!�S2וDhU����V�#b���2�M�>mWr~�,˓"���rOѹ��p�DK0;��0K��}�C�x~*� ��r6���uH�LL�i�ҳ!'k�dSK�c���A�׷��:uû℄{��������ӻ�	̞�J��/���o�j2L
��ڒnX�E%~5㱚��O�M_�"�q ���N�j�)����$�o=F	gO6F��-l��1=�9�b'���}H�8�N��(�U�7%)�����/�Aʊ���+9L�vQc�q�F��{b���Z�6��k�3d�^�����W/���Þ�ʄ �S�����~6
/�b䁂s��6n�[-��	�aU�<_g����ׄ�����FpM�l�7�+L��W)Rbǧ8�y��P��5o֒��[��e}���+Ѻ���0(L�}7T�#��a\��TlBu�����I��]����j���q�$���C��Y 䗄2è.e?��3��7��R�uF�~	S���>L~�����H|�I���.dy�.�c�Z
Ua��^���c������AU��$y���uUU/��ފ��?T˭��!��9`E�n�zؕͭvB������F�Օdzs ]��d���ʮznaF��<��ש�<V��;z���!�{���_�*O&������-�ғ�
f�`�=ʯ��r�'D|( }wi;qm�W=B*|��p����/�<E?����b��� ta4r���#dz2pZ��0���OqF�J���z��R�)��rC���1�/Η9�����u�a�V1�%����Z�ӊ�2���u��H5���)�'ԱӀ�#� tqn����.����<�m���jˌ<i�z̸� ������\�w=m>��� �ʎЁ���0�RI�&�ͫ$#��?edD�2��&²�L�2��{��&�G���v�D	r���m" ~�K^hQ�|�!�����2�	�ύ�ֿ����hgLҽ)v�SS0�ahz3L�!�u>-��ԸĮ����T�j�1�em��?Y�����R�]��ƣ���PL���0R�4�XǍ�����7�q���7i��Xj;����?��]�z��؟���p��`�9�+���0,=�W��%�0,XX�'}E�r�`�7�b��k��Fş�T�Xex�'�qrŜ�;|�*���ԗ�G@�Ds��܌��T���ASG
 =�HիXy�3	��}���ݷ��1F G�Z�����I@�܌�`R�x�7�޾�τ��� �4�;�pU����;&������i�����QeR�'y��X�Ե<Fͥ>&�[Uq��x^蝾��~^�nn�}��%<����B���Vʒ�r�yi���`��"5�J��	l�I���x���	�)�ъe�܆���ء��B�ɀ[l@	�L����Ӭ���;$]���>���8��b2`�G���o��֍ޤ~32�/�A���}�����x��O2��E��L�*�xg|����ߨJ���+��7��E���^I�%ҽ5�o���Өb�"��A'�f^F�E�Rw�M��C2����2٫����I+G��.oOq�H(�jꚃ�:�636�W��Sְ/���]W/ lgZ��"/�K�1�L�\�
�����É��#�'R��)<�\>5�0g���� o�\3;]U�����z��^#ͤ�O��4�K�̤Z�Uk+�g7Z/�;�Q@�Ǝ�DR�
ϔ��w�+��ۮ�����:Ɂb����?΄(t<���{a[�)�g��Uu� �$���#��XJ�V9��f;�:x���B�c���.�p�
#�٪ ��3���,�]���S�X�!$�{xO�����;��\�����ڙ>�,��(��SڜERT�](�C�N���h�I=��.�bFUw��S����+L{I?�z���
Q���0#�,��P_̌�f���-JoM�֟Ʊ-pX�0���G��T9}j�l���ކ��Z��f�V#���ޘޓ����`[-�A]7)���"� �sh�Z��w(��SZ�m&->V��*�����ǅ�FpL�(������p5�@�ۛe�����`?�~G6� 
]��4��1r�#=9Nv"���������c�G���:
��[���z�IY�` %O��Ƶ�v�pE�]������1�׽��4�`a�'��r�#�`�;~Q��{���V �Ǟ8O?�ȴ���H��|@A.��`�t�h��;T�3�����È
Љp �H<�^T^����i	��w=?$�L���cM4�\��r#��ˎ�#l�p�UG�g�����)�U{�_��żu��5y�e��� Zv������̕4�s8��K6�w��iGpoxԅi���/��+��V/������L���BW�>����)�`��Q��y�>�<G��{��p�.�(-/��}���G�j���_�`C�k9�1Է#����,�v��!'G��Ѩ!�]��U�|HSʔ�1��W������ഇ��]>��;��9+$�A'g1���e�}D9T��s/�#�]��;V�H�}mn�V���v���|�s|���������,PgĜ;�ha�>�9�k�S%�>w]Ǐ�V	��.��Y��kJ��|(��^7i�����r��W�Rʖ���m������J��P���9����Oln;��+��N(�sՌ��崵��yЉ��6�y�3��_`X|sX���Q�m"�� i��D�kͧ~��Ƃ���'3�7˝QG&KF��
��껪���0�A��Tf����wy|V�2�("�uC��[��e�n�R��x���#I�#�;5D�2��>U���.ɝ�`��$JϦ�2# x�`c�`f}�M� �O92,_\���"OGX�HXU�������5��@�)z�S&k�X̑����I/���e��i�N\��'>�-q��aR(P�+-�3J�,2�W� ���f��I4p+��!G��c;�%��?G��k*��Bm�bϚ���dZ��bܓ�%=��ǐ���Yq����}���kl-�r:1>�ǩ�����YU��"����ߢ��I��V��W�c�@/��X���wo5p-6Ѽ?ɬ��%E~ܻ���/���3D	m)�}��M�f��>&j�2�ˋ�O�.�=��|��&�؅B��,L����I>g2�?��Z���1)�\��i!)�ɞXE��2C�Ğc+ �r�ɻ����ؚ+�Y=9I6��RE�Y�j׾R	]�x@m�A�U��"|H���y��S]f�Aj��6-�f��(��ў�%R��Q���֗��K���UJPb5�К��Q��=��te��';[��FcÔ�uu�@�Q�E�K�M��F2O����:�R|���π���ۛ�H=����ͬ��0"�0�^x@��!Ľ��
�"��>ܼ2o�R	G��c�bC���&�����2)� �qGOaT/�O�9*��1��Y�%t�|[8��l���<{S-^��^{t���i`!,h��[����#5�nH��\�`&�����F+9��O{r_WS����_[iu����С��b�١c��kQV����?)��t,U�'2�n�Ő8�SD� �[���|�I6���
��(�M�2�_="Ix�˄fW���a����5���˥�﫯%��z��
*D�Y��3���:�V>_]��mཛ�sF� �_q@_�)9�~9y{<#���.>Ko�n�r�bڊ�7/�.d@2*AԿ��Չm�G��,u֮�Z�iS�ݢ-q�H�Q�M��X��J�����sE�i~��g8��+����ށ����jZV�kw���69�����ՌJ-z��Ԟ͟>vG4ec/�eⓇ���J�N��T��y�J"�- (j�ͯ�Q�
WU5�;%�in�]�I^��b�{�R2L�0���5H��GSZl�,��&�~�w�m'��'��^��Ԫ�BI����h,ai����7�M��[��L�>�����B��Pg���#ސNY��)��	+�·�2(���^g&�fxX�h���g/&@�1H�MOo��1ڬ��J�{��ݡ;���>ӝU�\�w��b���
��rEdOep,E����l�7 c�˕�<I2^���ʡ�I��#��0�v���_�wH/�wI�ti;�9���j�V ��{��R}�%.	hf�˺|@i�����K&*�+3Cr�
L�i��i �(*J��,�h��J
j�?�����ZC4�#_�1���D���f�7�+��d�����������qV�>��{f)#�o�@��N�ǵ��Vq�H�s)]��m��Z�����HzE��6�Q6o�N��lEY���*����c�"�#�X�vF��sHʠ�ؘ�����о�1½�Y���NDI$��	���� k#���u�+��o��֟������Wk`q����Bҿ~8S1�P,X����<ݙ$k����9��%�߯������pe�m!�����|�����mc��)\�����N�BN�.��ݤV���0�	���e	o�F���C�X~^�[�Mm��7��$E��
�qo���m(�S%3po������������㓰�-��S,���]�`��q�G�^,A�#ϫ&�;��DS�l��k��}�g��.�Qa�Z����	u%��FFBe��vp��P�� �������+t{�i$�L$����Cf�� "|��Pv�2 ��uУ���4�]K�=�����մR�M�)�+~�_�l�,�	+\-�Y$U�-���]x�jdVr�
�-��q`�E���G��(�%*�:gt���ie�9tՖm����G��D`tD6����S(�I�MA�tP�䦰m:���e/��R��R5��f��YXv%��X$�������j�7(���b���CЁi�CwJ���YB:h�E���_��ԕ�F��A�b�=�x�����������D�o`��2"h��C���{2^���U�06�~�W�\����0�Ѱ���=i}��ӕi��ԩ�(�x%����-ït��N�Ohv����n�O����Kֆ�'����^B2���B1�e��_`�{2�g.�s���NH#�����%�+�r����Ԕ-�����R���g)<ii�PU{�0T�/)�6BB��!�C���53���h�=�Se�m��<�~:������'_�2���$ u�#����F�d�w(�\�>3xɢ����״�㛹δPϫ���ݶ���!�k�u]��d�'#F�H���������HU��1�P�Ӳ�p��!�	IW2�a03��\E�L��/�W���G@In"�F�j���;#s����=$�ț�\#�����Q��_9�7���++��?�^�&�l����jN5C��;T��-n��.x�r&���Zr�5����?�\�-�E& �Q�����Ϛ�(��O�����PP�5y;��q�*
�MYO,#��4�-#&���T��"���~�����P�xo/�>��#�5�x��j�#�"t�"v�'����ű�����L�g�ǂ������mH[��
]C�ɜ�X
�H|�(0�cP�#_h=�E�ޯj���đT��0����6�T��#kM��UO>�X�)�G𨎔-�"G�=�;䔀���@'R�)�쭪m�^yg�+����[J+&#t4.l���E%o��mS<W�E�ྥ8�l���c��s�Wt�}��K�Z|�#����DP��[�'k�cH|"B�#��Í�F����za��}1�.Z�q5�O��[���������E#�\9Y�d-\ΙJ���pp8QÐH㹝͉g
�~ܚ��N7	�S�u�R��� �@����K<�B��~�6���LF�#Q�9�a�p Є��t}k����ڲądsU��'�eX��V���趂#i �1�$�c������5�ѱ��~8�:� "2@�� [�1܎g�B���J��{����s�c�R\�N?}���%��͓JeԪ��s+�F*�]LF�����{��⾿<Ipɣ����AБZ�r�]��\������ns.��#.� �+\�]ʈo~>���#�LH�j�;F���_
����������<��3��K�QR�뇽()2�_JG�[��"�s\L��&�3�4J��8���L����]HtU�=��߇�֝�v��?4&m��ǘ�o0���H��O���^��^�5e�%����dM��1���l�x��q*"�5���}�'	�$Ga&�3�����p��a�y�s�A��`R�\�����|�$�L�ɵ�R��Q��6s1��s������b��2V�����n(6�H������Fo��ϻ�3��z�_�\�4d���,��O})���f�@XOK��7T[�S踪Qb**�儠M�B���O�D��uV�_�[Pw��� #����S|�Bj����t�y�1�sc��t&šv:;��9�i �&.���=���Uŭ��#��#G�ѩ����Y;U�B� 	��4"y�&��x�5�:�)�A������\ٔ����fF���T��3 m>aZ��)�-�$F�/�1�}Ѳ��Җ��6
X/V�f{'}��K�&����K�9�b3KΈ��o��s#b1y�� Ob��W&UU�֨�>�oǌ�8���]L*_w��_~0�И�^!&V;�����D0q���`o��y͋�s9����r��&��f\5i� F=�H9f�E�$r��%v´�3ye� ������B�F�q���4д��r�vj��/�	�&�ja*����Ǡ'�$��}�W����s��-\%��N��Cà�ߚ��}}�a����@0u=沿[��ـ�5}���>/��!��J�������^)7���˛8x��f
��z#�~C�2�/�������3�\��v�%f�yԞ���� ʄ`#j7�����,:I�׵ZD�͠�}���m%'���:0]Ϝ���kl���i�������bJ#����#�r�*��(�`�!Ȳ�^���̉/L��ht� ���=M�@�I�U�'Uz�@�� 0��ay�����AF^��&f��乛�%��_m!�`I��(����e��=�^C�{��Q�a&�K*��Ŗg�$9�?_�t�m�y��"2��x�-�Zyk
���2F}�x����%�)U�\@Oӫ �@c��.b�r����1�'��ҕ�,��zp�>�j��$c�[��>��~�d�i�\�% I:��O-���|k���uh��tL|p�z��.Tۋ��$�Tx�`A*������6�f��~7'K�:� )�,������/N�"{�%�]��t~�GH�s��ۧ�p�jo}�I��wG�H��|UY���k����;7�HUn�ˣ�x���+gd��I��y�E�\���q$1@�򂢪de��F�f!�	:а.�7��G�$i�~_���]��8�6���� q��g���-�,/��kZ\4&g*(WBA��q����?2};���R�{���n7΋�PbX��˼j�d���S��/�ױh���sb�f8>�)nwh�[���������b�X�Q���Z� s�[�z��T��L���)�Z�Ƕ�U�;�R|Qr}Sp{ES�AD��vW7dPE��ucoH�U�.�jR�"m��~�����'�?7��M��
^�����ZJI��#�M~=��,�gy�4������s?�����1�I6�%�n`�8w�����i}ÛBR��sU�Y�D���Y�� wO̗��E�u#��4��`�_hIN�㣣z��.�n�֑�iGUJ�6��ޚ�>Af�hq�Uy��TF���ABX��f��%��B�[�;$�bV�3�I�Ke|�~�sJX���]D%��_��0�>����y�<^b����Q�.�n&τ"X����MK;��/��W�U����P�Ы2���^=K��ٖs!o�t
�p��?e�~d�7����}J���!ӀI�ꒀ�Pv�=|�7�'q��s��
����igƽ�D�<�.���� Z��B�|���k;�2E���+�x%76-�����?��d�(.�f�}��'j,=^�Ɵ�ę����XS��T_���&�':ڔ,y��*�ҵ��Y�IO�*G8K2�.��//��L*��8���B�C>>����un�J	�$s>�: ,^��!+W�ޒ_�`��DOV���@�˳�A�
4P��Az˯
��t�<Zl-��d� L`���>�&����ю�6�>4�hk:�kѹ�I!#	� Ƞ�~�wOG��Toђ�ȵ�ߚ���|]Ό8w �_J'�y؋Y�W����	Z�.r���P8�꿯:�I
�\ /���9J�4�/�U��^�\�>�E�3��(�F�F�X�_2/�Z�rv�P�@�� ����Q���9�hyZY��Cbn���B/�oc��\�:�<���M�O��2����V/PAdl�^�o~��	��~
�vz�m�M1.;���V��	@�$�����3qʏN��b��)�→m$���pO՛}������?�Od~F��s��!��U˕��ʇF���*�@�	D�5�L:�sm���<W�����^�):A�ӯO�n����"9
�<e����s�L98V*�QO�R�Os�F!�~�~�2˳������޾Pl���iA�[J�ޗ�q����f�sjSu>b��LE%v��<y�&?��K�n!D���`�4P`���~��h�S �}:���4BzG���o���Gl�a�Y��_�e?*U8�tǗ�H�rۻ��\Ƿ�$��u�q^	K��@�9;�6%�c>`�x�O�����'�oe5Ƚ��� K9n_��</�('��FֳA���N
Yw#Rm[,�w�AX�a���^ۨy�:��tU�e��+%�+˟C8Tǒf��b�����@"�uCDTQ/�pnB���S9�Zp��A�s���{aL8�|�-�����d,/n�{�IN�A�:�x,��lvV<j���g@=�Y�")s���j�j���1~�6&I��V�TcӀ���i�K$�d\[��ИpԴ�M�C,$(���n#�[Ȍ��~P��0n�t|ڈ����yQW%L]�J�uh<j���;����3e�WL㉟��|��%��X����� �<��)w%j䙦׎FV���҂�5�?��:��r�\��t��,F%���+���<x��坞G-n5��W����JJ��WO��a��R%  M������2�R�RSbc�8��g��VqVO���t�lwZc�"oR�<K���qQDyB�z�u�Q���>��>�n�e��A?�Կ�-����C�����t��/E����Cl7��]01��i��\D���%}|��]�{DxI^{���;�}���{���a�>��H�$�9#k�Z@�?�e���f�	�!x-5j+���X��m뇣���(+�,߅n4�E�/}+*�^:��[A�j��ʖ�z���������G�H7{?���ʍ��}������c�$�0�଍�\��澲�Frb�V*�[�VZ���X�JY���#ޅ������?�W���^�5������Na:�7^~�+����렯��i�w�@�$Z��@-�s��&s˹���eULO	4���CJ�N����o�6��(��Ϩ�:C�F��h��]�v@0�d�p: '\�A���}�&9r�)^���MVP�v�����ru�'�NA�qe`� (�>�?G����m�L��HU8b�f��r�Fy���[��ϊ͎��/-�w4�hM���2'��1��o������(��_;����X�{#-mL���I���v	��
A8
��ϵ���3�u�P���������*c�K�c�f^�r�n:8ܕ�C�N�̴8ff�V�{���qht3蹠<Ob�4Μ�>�O5s�A������B���?��L���)mQpi��:��u�$�'��8�v K˒걲k��7�~N�V�
 vPzXRנB�,���n~�~�$�0\E��DZ�crdȐя�"O��֍$R7g�X^����'AWF��$����&aR�����4��,��
1n��/���Z���{�3�m��
��D����Xк�z�d9
8x���v�"�����e禅y4�*.�s,�&�g�K�V]F�d��Le���@�ph+�Ֆ����*�"�d���Rl-����2��Q5���؅Q��Dl�2�c1*�|��_�bb/]�'$���t�@�s�����8@�l1��&�mh�38O�LO���V��MЎt��1��D��c����H�ϲ̮݉u�#�7�|��!�Ƞ���(�w,�;<�X�����j��^`�����>v��N�z��'�.Su[�0��OH��0�Ggi��(��d�r�~܇?� +L��#�V�_�в%շ��W�� �fi]@ɼ�[p��*lǔz����J�E�;�.o�%�|\>z�R�Cw-R�2�ʷ���`��"X��X��J�oq ����M��'�ne)��b���Y��?k!� ��)}.|�4�� ��<��Oi!�� �̧�=���'�Q��b²�n+Q�A�
�A0T�n?g��$L.Kh�1�*��uտ�W)\���T��#����q}��%jS������H֥����)]yUN��2�Ў�]�� �D�ޥ�Q<��ͺ�r����!W����w��0?�o�wڕ��_�+��|�io��xT�V��Y�s`��R�߬�`���	���w4���tK"RД��PGGn�0���k	#��S{ye��t���+�Y�0��F�V`n�b��ߺ�a�9�1�S��i��� �Q�gX���~�E;�0�i��i�����ʗ \��Q��wA~Z`�N���T
�?U�c�)�!'�Dgg(2�wH˖2/��.���7����3�v&��?�D[f��ŮH2��?�ĕR�-�	[����,�|�2>��[4��PC{��+���S��5A]�r��c�$D�3�M|$m���)��e�C1�0���|]��4�_F���A�4�(�Ã^�S����9��	��;�qu���.�!�T���lGM[�=6��	Jro�2Y�G�Q�WP�j�sL5�>�m�l��v�\v�<!Q��0KN.� ] Q����)W��/��,)�[z�����h|�h1�^p��4�%턈x p�hߐ��E|+P��/������q&��t��LQe���ĐĈhi�z���ks������R�6T��0�5L��yC���� y�y�� ���v,WQ(9�e;H绒"L[���[��#���'�}��;��v��i�R����'���ف;vTd_-�J.��*���8r�$�����H
k4D�=I�>������,�'� ׳�'Ƀ-M?���C�.Y�C@��|�ɧ�~pZ8���Mݤ��	��������D��O;^n��ހ�*)�j�p\IY��gv^&&]�������R�;�@�9�Kx�4kmzdY9kz���'�_ĸ����Nzxa25��^T� ����Kr�O{��l��<��0����u���_b�	 ���̈Ztɉ��ND�#{˄髵s�v![�!��̃�$Y��U�q� R��=�V2Ȓy�y�JZf��no�̝ôX�g3h��*	�S��3{C�Z7�8U���u*�t	���$b�bnt��. �5�6�C�'��Q����j�5��Ř3+�S�7�����V>A��X�j_���ۿ/(���.��?�#���aV�8���a��C��ӿtU�D�W����X�v�YUC��=(�+[�L$�$��H�('�>�<vك}sf��qe���KP ԉ\eO���C'h:7�;�F�䦃z^p���)����'$�<v��A�F��J�?ɡ'��ӫ�	Ⓓ�<��(�G*�H���G(�w5�2�"��i=���y?���͹j1��l4z�(�Y~PY�yo���)wh>�E��7�h�b��c�1)l)�����a�}����M�O ~y뒺U;��J۾S/�w��X*��ߕ^�>u���l��k`�`v���Y�~<�R��_��~h����9��C����PJ6O|�����߆/!O��P��}�|*��I���G�B�������
�{0�����,T'��<i���Lh��^����qW_�s+(@:�u����YD�:ɐ��n�V��p��7�V�uO�{[���mW5Ѵ���ܻ���P��o�Џe>g-䣍݇Ӫ~#Ӡ}��V�Y,r����-�sL* D������1�5v �i0�th��䷭Α3
������z�~|�V}��24�^�y����Jy�l̓�A��C�)���B*)�n���RcG�&����$t�NFgD?~��->�)�� /��d���?peԗ���.4b�y�\;�W�X��/��ۓE��rtz8"�:�~�lÓD�ē�赋z�Y��ޑƜ�Q���_���k�6B��DqvK!��*[O ����˕;M��W) �� �#��W�vec&�VX�q�d�$۠N��� u�J�	C���{}݈�c����3?��oX���O������\Z���F��VqZ6\e����l��E	{|��}�y3G�`|��3�]���V�����+��	F����;ف8�h08������s����lFRl������i�T:�o��/��K�=-{�
���O���Y�qo�e�E9�.��d����O'�@����D�� 
���}an��+��wr���%��եڭ����)og���+�y�H'�Pc_��|��
t���`S��?�N�;ՁR^��~W�ֆ��B2G�NK{=I���9Jd%��/5f�<,:J e�+Lov�%w��L�ACjhMY��p���vx���>c}R՗^��ʭO�>��	�t�f��s߮�~��#RZ�Q,�$��Ť��r��Ä�l��òR8��cC쯦��G��c��K�<c8B���}֑�AO�k�:����mZ7��*}�L2�K��bD�;�AWP�Y�jL�dE�h�[|���CЊ� ��r������b�Fj�
C�� D��p�3a�o�����a,���Ύ��Z���P.M!���W ־,�T|&�=�0�$++1×؄��t|����xpr�g� ������H�U<��">��<U��1�X��sۆ�֏�	�� t��H%Y�#��m�񠡇��b�z�ẙ"bj�j���}���0�i�/ G �?	�s�rY`�O�=��JXk��
�"U��~2��!=��-�3 �1u�6_�w���7ޢ��&�����m�Z�r���_Py�w
�{�n�g+`��`5�l�N�Q+���Ó��fu��ڢp���ti�F1ѓ�_���K)���<+S�ɩ�21�o6���� ZRެi�)�H�K��v��Ů���J���`��	���0iq!��~��ſ�"n��N�ݸ��G�'`�BwP+>[��c{�Y�Sos�;��Nk�2�(��1����Hۺ��DiO����(�"�q��t���3d_�>#���bgd�Ѷ�0��R�m��f�9L�W��sTWG\���G�)�u\O�;��7mLỦڀ�z�!�_R��}ܦ�R탸DJj�cN��^	8 E����>�^�O�<�6�!�k��JC8_�o��;Xh����xo��~B^�&WBٱ��s]�3�<����f��y��+�����C,K~ҽB�Q
���� ��.��p�'���B*k�ӥ� ��� ��wV�W���`�G�������n��.u�"�_�S|����Fp������{��99�t)�&�z@-W�w�k�����d"�z�7�K�!I@��ba�yZ��NE¤Ȼ�]�G�+I�9?6	4����g�Y��U�p��<?y��<�_�5bz%=��^|P��e���?\M�z�_��̂�@ب�@S_U�^4C q�(�D+&>����I<1��V�;��P�P�/M�����0`>��pl���F�r@i�����oM�n��_�V��b@9fmX<S�vRE�-���l:��-�AZ�dϙ_���}"�\�`Z��s��ʴ��m����EO�|�s�����h��rؓ�}R�2���!�#�So/?�|����d�}�:�9����gED�3��:��x��M�y���jD�q�0�-;rλo�D�d��L	�{H<
���$��+�}wr"]H]T�Idp�Mm���n���|�a��Ap���b���T�a�l����\I"��ǰ��3�i��c,�yL���6v."�6��B(�;z����	>n����b|��0Au���9$3����PU���ea��RO����և|^�16�J��FE�E�p�Ye
�$��7���!���H]���H�|G�� zU��T*���ջ��P����/�)���sj�>ҷ:�>���5.��X�*<(�Y�%x-;�n�<��+�=@k�N+I�BKK��&o[\�'�/���-���sV���1��pj����s�������d�$֬�p.p�H�dꪂ+�UT�x��J�$�|��gA*�`�:��Q��
��]�h�%&p�vq����N�j"&1����v�	c9\�MC��0uCWxcx��ʺs�.T�oT����8^s:$eP3���G�y�?j�B�H�Y1
*M�A�Sr��J|��1fr��,�wL�sO0���H���v���+C�����nN��֨u��|Q[�sPk�=�B���`"�j|0M׻m�~q�Zh~OD�t�ϑ�K�V��1�����P�o��K�c�t7N+�i��R_�H��eg��鵩��+k�p�e{�
T����Ğ���D�'�t2�]K���<`��𽖽k�f�P	�`ɨ6��p{��Ⱦe�����?��@U�ǩ�
���I�-�֖v^�p���s_�l/2wH잮z��m�('�o6��P!�|Z~�y�Ĉ�k:
��ٰ|���w����ƬR��<�5پ�6.��7�]�˸A��דf�?�3�� cݦ@��T�Y|m]4�Y�z�oO��-�=��+��ǫ[6v���{��8�Ѷ�#����B ��w�ճ��5&��B��C-� �������v��5W}���Y�L��j�Lt޺��p'����*h��N�چP�EL�V�k����,g�	Z�M ���A��}BXc����-z�_'L@`�jODkس���ƬV����I�D
�Y(��6�oj�5�%B��X�` �-˽��`^Uw�.������G6���~�sASw��X���<g�Ͱ��/R�^l�/R����
a���9D/xV\����VaG鉗���nmu\��UR�y~%�|�F.��$�)���hB#*h8[5|;�ٴ��R�y���w�H{S��I75�4�B�O�X}{�H�ύZʊ�_���d�;$|�Ncެ��;�,��;2H�q��zIZ��4��݁�)bvȟ���A�	u���q{����rі{���p�����c[�������6�`Z�@u��:Vfo�4�-���]�<�jC�E����[��%�V�ɷ��M�.%�0T�����u�b6�MJΙ����B8���{��Њ�X���=�F��1p_��ɋ�N�ϼ���eюlY����Zv�ڜ�Y���Jj�9E<�����~��ҁ� /cr��G�ɗ<z�]p�3�����6�ET�2H�9�r��fbQH�(a�Ō��$�E����^�C��qZ����D�J�rw�s���\�*�aN�PM�,�ʨ��26�0<����H�!b.5ư����j���=�
�ھx�0�<RAY��bQ���j8A����l.ھ�b���n�E��iT5A
 �]�C�2��#[�	��kL��V�̷���t�~~�0ljC.�g��b�@�����v�V{�*
�����]�]�y﬽5䟧�Pp´^^��\�����gT���C�3D6BR���b2����NG���,���u�� �ר��d�i� w���֌�.i�����y�"���-_�L�G#$������ٙ���'Ƌ�ൈ<�%F��:�R��Y�]���̲�z� �h��1�%̮�-�x��9�9?��!�ӖB�
�Q�����S�u
���|a�=_�bq��u���)�#zT�KIB�r�rKs_x'7zL���IGq`�v�]�v���p_���;æ�/�OΗ�V���%���S�Y��w;�����?�w����T��|5�e���Ʉ���x<~�e�L��"�_ƎE�sT0���/aqWz���1�-�4ЬY�2���`����0�7��8�����i'n�%.ؚ[!�'�QG_��N9�/��Q�hw�q���To'��(�ɏ�	���{VS�{B��A�{C�b���c���oħ����-(P����HB]@����Zc�����V��Y]��)Η��3T���1��~q���B-��Q�]F1H�l������_!���;����h��tL�Z��T�����&}�壒�=��4 x��M������y�{ܢrEP�3��ɤ�������>���ЭʎXȯW1�s[J��[hb�wH֑^��)[05E�
���Xv>�HÕ�R�2�eq�b�(�U��E�ƘQ���f$�S�4���fP9u�}�����E�&(��ǔqU�t�[-�f�+��A����+�pD^���_?^Tg{	�)u��Ī�r�=f���Î�8��K�����|��?)�o���1�24���2JW9�O��t��s���-��� �Y0���7=����4�6�~��(;��9P{g�0���k%�ʯ%���3�t��%{��s�|�~��a2B���p�_#l'�� �*/�O��Ju5v�z��W�����-R�0���T調ಪy�� �w�����f�+�KU@9�~ �h}j��������bwbR�SVHGl6����ő��q�_�rJ��6�sR+	�͹��g)��|��]_�ƻ1B}|�<���׍Y:�V_�Cr�UW颇���<k:mup��or�����[M���Q�P��o.ēe��{�D��H�ѯl�ֲeZ�Z=������s���� +c'+Yl%��[�L��7FHr��a�#KnC���H�\?�V�{��5�� ᓉ���#�W�z�  �
�����hc�<�����H�n�ʂ,՚7���+{U=��:
�4�"�?!- �R�e��A?�ti�|*�K��!O���>�&˵�#�]�)w=,'��g6a�Ξg����9�#����W!��w{�@^!(ze�{J�5ie�ȩe��H�JG[�w��HwlIw�P!��)��U�VFO�u�7u%�xM�
J���Ό�;a����֊a�v�#���/�N �3�o'�x��{V�8^L�B{����KD/ʒ2����;�
��ΐ��/��?�oęEV
�󋴕0�j��[�����G%a5��:�������D�Ug1�|ț�'��VU`oVփr�B9-�KI��N%hu.+ӊ��B-E��a3�|��@?��ΒeJ"��H��G�C*��I�_'�`" ����n<hf�} ��e'/U`o��P�E����
��B%ȋ�
)<8n�I��Yޟ���?�~"��\c����/D�<�ݤ_j/��D^�S��A��Nx��^��� "�'-��g�	���(&Q+"S��g�tj��S�uQ��n���ߺS}���5�4�JTh�v]5LOz�E��ԶK�c� 0抲��7y��RR�]ǷU�*�3.�p�t�1Y�4}�|.���mU5*M��t�NWU)��C$B�-�¨��g�[�4���%	���~���?�,�]jM����~%�!�8��#Y���&k��0�U��h[Kh}��m�(�"�����k_j�#ڻN1��ӳ�BTIkp
2ٴ��l�fȫ��Ƚ��d�A������JȬ���Ϳ)<��m��������)�&|k���ܥ��~�M_x��ց$_M�O �Y]��4����]k�s��,�M�W�P��m`u�V0[����>v�u�5�4�<��`������K�� �קT��{�]r��1��܋yE�A��-�9�����<�:#@�q����L�M�u�&���6Lb
u�-#���h��(Ǿ��e]�w�2�����4E�*m���]O'cY4���4�kw���C�D$o=K�f�
�ZM(B�z����i�6�lg��xsN��zN��c���E}��ҁS�k����C������Gr�S[��߮�"�Xn�'�)�:��]#c> /�m{:�1�%F��M��rӏ�!HS���w�B�$�\p�]BD���1��]���#5<[��$:>�aGY��Lk~���h�
��`�G��,mѳ'�FH��[�yF��Z��޷�9�*�����.,���N`�g73T1�s0`� H؃����������b����-� ���&�e��:���=��X�L��H�\��H�<�4@�!�%���+�I�ͪ=���F~�C=��z\Ȃ%�Ҩ� ��ƣXVu�{��.6)iA��E��!�$�Ͽ��wU���u$C3�:��`龩d������Ւ��O�+^װF/�>�/���S5���-��1*y�cB�O�aN���k@Q,�����T�8�Ή���`����G�)@�x�g�phB�6�����U+�u�λ{��I�W׶�Z�]�4�Ms���}���9����ދoM�`?N����)��	ol���P��R���zi�ó�d"�F������|U��;!���gj$�&���q)�.o��͆+-��Ia����Tu��
(�E5>�+ �����u%~H��
�R.�"y@c���I�P��B&�/�H��|c��� *�Ⴀ�΂�DHv��G���I�M���D]0���/�K��"|s�,�Փ����]Ka�`��D<�g���͠�? �4 ��u��7��ڼ��ok��.��Eْ�}���u�:�첝LO���I�=#Ni(n��?'."rS��a��h<ں��ձ�U��+����ܒA"_�r&<�)��2*��h|���迯R�<m�p�{e�(j.�N�n��;���%bBd��Р�<���E�;���!��sT��ߦ�'� J�T�R8j݀�ܬݏ��7N����qY�۸��
i�@��m������TH��̼!�h	V�����Q�ż�sϵ$�+r��������`sf����Lr4͊��H �1�����SG�O ��d���?^Vr�;�ه���&��
���$���幟�aE�>�JR�^`d~�`.�l�A<�0��u���#��T�[��Uyh��c���>�YR"՗
�y�5�F|�]�1J8��dk
M��?��	� `P���z�k3c���k>�@?Bts�/w7�:$��*���'��q�ۈ	 2�����EX��w��+�ZU=�kT#��3�^;�$$�P��֠��L�~H=�������j�L�R2Z���?��2h�l����6�.��� ?;��/��wȳ��q��;�s�f���p ҷ��/��O���;�q�=SfE ���jLY��8CeW�9�P�MtÀ�<gl-���;P��ü9.�3�=8X��݂�B4�����άݶ�7�������h�a���p3��BkG�I���*����a��§��'�>�����lg|Z�}�x�;��v�G(.%9�V;�䴯A�����(+N�p�.TB�O4fG�pC`��l������y_���
ଡ଼R�?�!�D�OI�P�,>�0���7�P������'����ln��x�-@τ
��W�yk5����\�����I"��P&��jh�H��G������e
R u�|Qȱ-���|����D8_ �B�z\j��\��8SJ����8�˹�i"L_�YR�-�P�k޽+AB��"����1�N�mf^m.��\�$��ˀ�<ω8� ��
�e�݆P���ƁΐaHՂ��+d�=2k���"�KI��wX�盛y��cX^J'��N[r�_�L�y��ߖ�	���l��=��q8#�SV������[����)����۱�N��n�_��Ι��2�zV��Yv���s�)��x[�m����:�FN��F�g4]�\4`Z�+�L96�������(п��O=�pF!GT1���)�e#�^�$Q�O�ʞYN��02/��6��I_x��=�˚W��S�O_$#kC���ۛ��VH�k_��y�����/�	խ!�lRt-[�硏/�P٨��lF`p'��{
�r�o�G�J
i�k8�T~Ncfڒ}�R�k �����;8|�a9�����&n��H�쮰5\*��TbO�LԜy[i\r�.���v�ĹIǢo��:5�i)˱:og�͝-&˩�@iozd������m{8\�״������ݫ�W*��-h��+a.���l��s.�F_t��8��.wj��P�o_D��7�3#c�D�2�y�&,O���_��,$r��T/+-!���G�)�n���6�v�qGiޖ{�|��P���h�����E�u"y�ѡ�*#�Z5^�*�{j�����>�ԍ�O��ϑ'�{�����)��J�����ٯ��; �j��Vi��
n!4�oİ��K����bI�Zi����h�E�
�/�*�!�.��O]2���q`�~/Dgn�(:w��Rˋ˾�7�������q;#~`"��F5
 e��o6_�:Jѯ��߂��U��-q#ĥ6�6�p\M���I��@?���f;տ+!L��8�L	=`KΠ��y+��jjK�Mk��+�����́����h�x��=/A,�OU�"o����������Lr׫��4���UtK��c#=�5�b���.�H���˻�K�q�����c�N�m��6�E�	���&�
ibQ��پ�L�a��*�G�3��)^��:ڹ��dLG��ej�VPr ��HB{?&#,P�:K��e����/~i-Zp��{��L2 ��U�w�P V���J�~�=h���F�,&�$�?
���	pƴ�"� ���"S,j��MnU�f$�Z��zf�<6~N�)�Ia�`�͝�����F����%aD_E?��V�$�l�;KK�-�4���)0���ŕ�ǵ10؟���8��K��uIJ�)�K����9Z6��>	<Ʌ'tP%�(KS�Ȭ�((2�z��3J��1g�6x:��ࠂU�f���T%Kl��=����Oƞ�Ǥ��S�J�1-�:���L�����23��IL�.$E@�YH��%:��(�����S^:��,U���YE�uI��%�+�z���k�w����-��]іL�G>o
��9�T���У�^w�r.N��W~�#�ώ�-���}R�JO�l�Z�PW�4�Ġ��ְh�`+1M�*xX���]��j�0*-K[�T��lkYQ���´�RPMwx	�l�w�&p�6k�z��}Q�W���}Dv�޳R��$���dw[7�CH�ҕFQO�����O��^z�0ҚW�H�jc�����8Q�(�
@ZoR�1i�gN�[�����}-	�˂k��/1ZC�Yc��&�;��z�}��2�Jw0�����1�4IK^$Es�@��"4B�:���y�����g�&��[Mr�w�{H��,��o�9�U�EX��s���F;���%��C��2)��CO=~�OU
�i���?퀼
�2e)_�!���z��(`��9��  �RB�[J��FXZ��;ϫ��* 	�)u� �c;^��E|��q6m�7�H����8N��p�"�C����c�|-��l��/�`�H��S}���2=�����P{0!�BD	��<���MO�;3�flַ%��EMC�HH!u�{)ڊ7���n�ԫ�N�/����aS8�ݞ�;t96�1����H�d�9�T����6�-�ȱ7�sRP`�D���%� �˰��qU_�+�q�q.u��JHB�(�<�
�S&2������������h���\r��x�*;��98�<�k�s]MTuCf{~����]';�N/l)켖Nh�ʫWo/�q�.]�ꮖHm�-kԨ�D�U�LJ�O*�.H+��5#g�݉�Q�,?�jpޏV��Yӕv���L ��#�~"��|wf�8dm�}	Mo��F�,O�ܼIƫ͜zx�5V������lB�Ւ��B/*;��M]�|��'�-dkv#��:�g<�<���π��%JǨk��}ψ��[MV�0��o�?����߉���j�$�H�g&:j���l�X��6�P�>���R�����h��i'��e{��c�b����,�E ���o׏Qy�a:bWN`��%h��H�S~�ď#�X���"��:�r�n�I���V:OG��P������K\pҷAD�:�-�%�-����J\���[�H�6�	����K�4e��(��b����6�#��v'�i^��̜^�B�f��Lҧbo��d�1��koa�t�(;;���Xd7�W�.�9D��IH��,���(�s]����k�WfE]ypVt;ԭ�����|�DN���~�>�j�m8��k��gb�����k�pL 	�CKa�����!ƌ6�/I$�5�դ@G�ӱ��mHw�W`�n)�b;�FY*j�@����`��r�zU�kUO�\*ع�	�f���5v��M�S�3Isd/�H#���%�6 y���*i(���a��_1�U�x]P�"K�:7%�k
s�� �w�[�bI�k��J��)w
�T��(%7|���ӓ��sbA�h��A���v��Yho�|��z1�3o��O�i'	�hfSy#�gPN$��J���pS���%�]��}��ȗ�B���������j���֋n��2k�ǋ%�㽑.>Ɂ�{{,q�笒���)����2'�2�?O[x�<� #T�(B�K2�}��ب���s5�����Q5�"��L�E�J[�K�Q(�PʢO�{!���� ׾�����=	Tk�3��`E֎#���
G00��4�1>�E��A�ߓ�7�̐�z��U�З�@i(J�$g��[�B���l���0�R�8+�GZ���,��<�`��r��K�ڶ�D\����tRԎ�p�=���Ng�Ӻ�
A\��
��Ws�Y�݆����m�O7�'�����&�Ї�	m�mْ��A?��z/�h��z�$�ʨ��"��/i��w�,�%:��Ƅ呤�E���,�.�	fN�;��x,+Ԉ�ҚU3{�[vH���%X^ȑ�������)6� ���MVh���R�54�꫽�K�#��?�]�8$H��_�ʊ|&��RVt�UK�'hAJ��
�J�L��"E�o�0�𙏤I�����<6!�,Đ���O^g�N:�K�4F�ϲWqz�J�u_ů��ܜ�1�4U#(c�#9ک�tJ̱Lm[�R(%j�v��2�WJ��P�A���36�x6�@��Xg��BG0��B��P�ԉ]�B`�a�&�ֺ$\f�fKt�+ۉґQ�J�eF-+�T�0�4�����D��U����罫{��p���O���oӴ�a���IT�|�p�Fc�6t�2�qx\�iZ��@������i��qL7%9	ZT
�P)�LNT��1��q���x�FӐ�f�s�E"�yx���%�3�15j���H��
��m]Zq�
-�� ��jRѨ�Cҳ��v�TM�	C�$ػm����������cez���cA�L�MZ����$�āM�D�����6gL�A��Q��m�R0�i!�Wg	��L��܎��l3<dՂ�ÌU�U'jf��ɳ<���5�O��Z3޸A�YX��ԕ��v4s��}��`�E���@?�����lU*����p���#���2&G6>�R�r�k1pv�t%˰�>
�D`K�jF�j�՚T��R`&���/|��6|��������SPٻ�p�n�.U��X���>n��2�Yt��j����ΰ%$q�f���>T)��er�w��Z�^��m@�[�[w�y!�.
M�͇�LG��8<Z��2o/��l�k��^���5Wx��/��m]�S<�ߩc[�×<�s��T�"�W!iR)��z��n!*�ug���Kf�#@W(|�cQ?�s��&�okW�b?1�v<�G�z	�%V�~�6oOA������ܨ����jO�
*8H�->�q���OM�_�T;��e���	p�=#�eS��]у~���U��`v�y��׀�Y���{K�Bm�`�
 xT�jp��� @gܥ���޷K�k���fa�����
�&A6����#�֓8� F�T#E)�:�u3M?��]�0�bin�l��Um��1w�~N�n�l����f�`�{�F�`�u)C�\���l�SD���Z�+ZY�jBU��f�7vFWuĸ<AP�(q���g7'��F��ݥ����؍�j<����]]F��42?��eP@�v�&MycƇO����e��X��4ti~R�p �CaK�"�n2�����q-�2���\/u9T�j�x|��A�*	�/����8j�����z�a�G�������"�$۝�T~��F'�>�%$��Ь6�O�Prr6*��M��$f'k�+4P��P��D��'���ژ�oQa�ٳG��x;<2o̔��4�d(T1��&}���P;��M���8��������5�L7R��
��}�!mPjپ4Y��_��K��A�"�G��<�C|	%px;��ye���<Z��0n ��PV����"1A�-/��m��V�G���&i\��N�xi%932.�i*~��)��'ڥVe�j����n��#g�6�v�n �����~T�����Q)���W����l���S�j��w�W�<����-�:0�P�חP�)߰�M1�1����e��@�͹�'��J[� Ȟ���F�n���",>	Л�eԉ\uhB�vPȒh���
q����3�p����e��n���5�{Ns�pL��B
�vR-�렔��/s[n��:תG�6��7e�?����`�)�@'�ü!Z�cU�»�� �2�iF��gō��y=5ْ�LC��s�����`�i�r���d��+[�Z�"F�<3�k�s��|s�,�s1z���.����]�md�}8�$	hQ`�H.�4#��` 85���f����u����� �)lZ�W��Td6m=-H�_j�6��n��Kc�>��W��ޛ�������9��Y�A;��g��7��e���ߢw@�>&U:3k���u ��*�f̻�x�ml^�.w��9�O�Q��nX����~�7������׬�C]`�^��v�k���u����~�_<6�#��NU�a���*��M���4/�o�D��6����ʖ�MT���@'@>^��P�p]]��`�دeW�C�PƎW�ڮ ˸v�/�ϙ�A��,}��ϟ�χ�%��nӖ{�lo�!�7�Cl�������5�b�xc1hZsT��Z8,q�-��(��5} ry���e[S����;�rC5ݫ/	ꡂI�+�Ϭ�#G���:��f0<�����z��d�j=�}���� ��@�=̽�'��`G�|�"}rI�dI�Abf�6�h��:�+��م=uȖruJ�n�p,�CԯS�\)����>�Jit�����^b�!���6�v ���[f����7|{��˰�������k|�e��j)�P�PL�r��lf7P[di�;p��".e�~t�
O�����h ��r�y["-Hm��I5/d��<���1�I�DO�,����/j/[�}g_�X|n���[V0�BZw�`�9���t�yu��d�a��+�:LGׄ�(	��
�-��h��G<������u��8�ՙ��ɇ�2�	�X�Lި��}M�|��?�閘�$Cx�g׺�֨�z�3�.�V��JnI!�~��Ṷ�+��EI�K���@��a��ZR�F3]���SN]]@�oۣ䑬V����~� u��7�l��u�����Tm�Z)!*�&�Y����K���Q������N��nv ��׿���������'��a����c�h�O�Tr%���	����c/f��V]��XS��IuV�� �j[�)_��_4u�B�2G:1ԃ]̌�!�y�ͫ�{��N����?#ƞ�EI3�V��p}�i�,�3O�4A��;�{�%�X���?uʾ�ƄA�]d���~kRn���Gz~~���O}ֈa�Eػ�&�Jm�����*��������e)._4�k-Z~"���R���R�er��")]��/�g�������>�Y���
��Л�͋���v���ńe�6@�=q��-y�0��a��E��GJ&��/l�܊0�q�>Ҡ	��0�2�]�t��(��zy9q��>V����9O�n�_��|�fJe�ԽA5
!t޽�T����G�K�V\���{Y����P�$��1.z?�Mٴcs�g���T%|@�D��5�j�Nm�Ź�$(�j�����>�K����Z_PP���)��I]��EŖT��[�7��sPtY*�Ҕ���$�6��yq�.�bv�Ā��[���7W�8�p�Qɣ�h3�hF�b>��TnG��%�c��we4���ͳ��=1�����tq���4JX2߻wA_"���-�W-E��~�"9���*���1�tnn�ll��c((�}K�X�E�:���_�b��e$��e���0)�0Fѫ�>
ν���фb�[X@�����_��}�$�F�Q�/W]��ZN!���_{w�N�:Y �Ո����+�D%�h}GX㞒S����=ʲ��Ɂ�C�mn:{�H�������Hzw�غإ���_v<d�<\��V��81N�SmZ�O�j#���n r�`�Km��u�����z�k�lӁT�bɄ����Pzլ�q�%"�ka�}<���mw!��Mٰ�	5��4k�����7����!���Iog�W(��� ��0�޴���E^Z��ПC;!�֕�K
g^�0��^�A(��U���י����Hy�{��n;��5�7�P���`�f��#_�ƈ8���O�Y�qn�#�2��5!kt6~��b4@�Ѷ�\��4�z<!>��U{�}�	�+g��SԊ�i?�E�"Ǽ%�������Q+�J��(j;�|�b��B�z�tc��y5Ke����4���91	�{"��%�����NN�F��R���s�v�:��/�6�k���;���p�s5�78�"IX����@Ro{+C� (�d�k��נ�(˽�����Ƈo\��z����k�꺳���˛ו �݊�B,#u}�;�}{ٲ�(fyx �%U���y���w3c��r�eݞ�V�����5d��ʭ���G�X	NH���e����s��Ł�Cܷ�A�o�WY�g�O�Ux�t�n�x��W1��jhv��<��N��*l��c1�=`-�{����6hbx�.s'��C��cR�������<G�B.��`H}��`�S�`�����hO!�~bᐫ��>�%��v�J�f.��*�!��<�
^"�eGk&��D&
EW�~�uu=x`Ɛb��9@�̑��ߥO�e���˅��Z���S�����ūG�L��Ѿ�'�<�O'����?���2E�o*���r����H��# I��A�_QS���J�ң-�q���k3�i���ouP��ҪKXe�*�ry�O�f��u����DB�'l���;����}�KN�����8�#
L\��|L�uK/0�,��󚄋�+KؙÏN�اf�+d�u��¿R�B�j��S鶉s�S�hao���L��w��q=�Џ��[+����ٵ�\jy������`�mH(�U�=K[�вn~��iS�N���o�U�&��_��\�)3��@|��1�Y�r<�;��&(h��O�	�U�lvS�ޅ�j%_4X��G8{LИ2�?����$��T�+���V>r����!\̌�0�6I�#*�2���E:"R�[��|�ga���o���T�0�ŭ��!:�k�kB�\���D�t��B���L (���qM��4��f��

������?�l�����3��VE�L)��*I ڢ�]��'�╋A��6��]��}"R����nv���I��n"��?m���5���q$o�x��_�.h������7�'߂8gF�+W-��N>����\�F��5� �]���pxk�6,bK��}I�85��F]8�ӷjE��ˉ��O5�e�k	���D-`~8�I�쀗��rM�ǚ?bo8p�&N]������]SX������L�8a�]*�9���E��!n���V+2}�j�L õ���ؽ�{� 8ƄeY/�T<���4�#���49~Rk1^g��������oa���h5\�9!�V'+1n��x�2�t��p�/���NO����ݗs�-�TV��]
yL�G��!����mZ���>8�W$u�1�����x*E�H�	XS��xAj����N��E&��{Y��:�\b(���'>N�]�3k��.�0�hҡ�pTn��V���o@]<?+4�م,v!��T��S�n_jv�%�����՜l�h�7��By�U����!�M�} 2'��'���	�Zh��U�5�g�����՟�N�
��� V���:��״���`��= �[s���WU2,�m���=�l�c]�1��p-	�M+!2g	x�e�E�f_�I��R�|%O5v� O�G[QٯJ�?L^~��؋W���WT�\y�w��HϚ��FK�۞w:��UD��V�Q�<�f�+n� ���<��m���ɍ.N����!ٕ͝�i#��]
���wQ�Շϗԗ��=!�挍!�$d&�8�Lc��`	F�> �B�%N/�>��:�q�#E��A.�/��F'�wo���/��#���{�8��N�Qݤ��ج��}��u�5"����m�MS����V��M�bT�J�2���T@�gܩ��%J��n&� mOz�ɫ�?�ZZ�T��ֽ��3�-�iM��z�x��I&\~b:(?��놸!{*�p̮�I%��B�Z*�y������������BlcL�G�v	,�%��ћoN� ���q��NQP��-f86�k�?#G�c����T�n�l_�˷>��-4*���*�����my�ᒯn�����ك"V��t<��h��'�}/��B��Y���&�~��ӧNk�/�1`������JC1�#X��XI�.�=j�~G��������RU��Ye"D�Tk9\� �y�NŃ�F�*�(���.��+��-PX�1,�Y�P�SӤ�6N��}�O�S맴���J�F�!+$_���rd�zNg���:����33�����j{y��^�$�$k�)@��_�=��?XBZ._δ<�C���1�y5��A�����&T�W���Y]���m���R}�x�81r��%�&�"?]jTOi8������<D��p�	��ל�w��=>v��M�6��M�]}�B����� ���u=Xc�ZO�Q6J��'mF�$]+e��]���(V���B<���kV���)h��51��FG����������4'�9�e��_���S�L��؊Bϛ���!u��/0�-T��=G^̈SH]k!m�7(Cۦ��"mO�mC�#7��k��󽸄;�"M`����
��ނ�.��QL���}tփ�#f���8��q�&�]��Z�� ��!��B?�!��T//jE�A�?H�?�P
rP�dY��?^�1Gٸ����_�d��<�{��ǐn������B����$Oa3�G�ش��V��s��b;�ݦ��$y3��:�d�	��?Ҝ�r���.Ġ��Q�G���AV�v�pg����桞�J��o�RVU��D޿�F�����Ts(�1:��]D�;jp1��"3Z��b���|���H�w^���jQ���L���ox�;��:O$j:�Y������KTX��N�c��Y�7��_�0.C�e���
��ۃ�'��-����6��c��!i{�:Vk�WZ�	}�ו�n�(�8���ɣ�o[w�������.8q)�4Ӊ�l("]��d"��?Ľ�>&<;�O��.`u�o�6�Qi~��ui�&�u�'p�P��#�#�H�F8#����e�AڸQ���I^�C��+┄�/���K��f�"Ba����d�>��p1��C ^̤}}Pn��ʵ����3|gE��Ӎ��K�z_M�W.�b�jK�Ƒ�;>$�y�M�D5ٵ���U��kxވ3�#�����@D]�9�ihKC&����Ď$bz��~#j���{�H4$��=&(7����'��M���2~nD��ӑ�Z�K �L��dmC���r��C��q�+4,�P��غ	D����b%H���7��D�|h76@և��w��s2��Y �U�+��}d��"&�!K����������G�E+"	t"x�,�&xL��o*�G�����D-F.���Vԗ��%;ΐ6T$1��hq�wJ#Rua|�m�bLs&�} �Z�:��F�u���� �������)WB��mi��z%�g*�8S`<=������"��
jB���������mB�g�[���r�Ɯ�	���S����u��0��[�~�c0)IA_�uI�&!]ז��N��[��x��eFŌ�3��t��M�A����_�ϳ���K����|������h������3�i��+�m��>p%MY��S���F�)  uYs��@v�����i�^�B kMy���\`��?�}��zWu��U�k��C8י���Pu(��&(�'�,o�V�Z���$�X��_�Lq�mc���ɷ�{F=��:�1�chG|��T��ΣՍZ�S�\X'�T'�}���Z�/�H(u.��OG!�f��}b����U�Խ'f�>B�-32����1'Y���I��Fwܱ���&A���p��^WÑm��K/j���+��_��d��g|�M�f��8�Y��t� i\�Z���� ~K奵2��|�xXt��y[��-��( ���%1'�u5�N/����L�]L�v]T�7�i��DXH�3��\�t<�;n�Rs~J�2Yn�%��p6�>�4�xi�0x O�H<�Y���R�ȿ|���[.�c#��6����Mi�`;�Fؙ^�F�8�`Z�������u��1m�ybe_w���cǿ;f{��[�	��<�fS�$��|��? J:ONv�,��؎]��DVVz�1Hu�|O��u��R�Յ��{ݪ,���K�2���t��w���S��E�7�F�u��jk�D �S�����Q.���m'�]Q{�n�0��D[���o\H����(:u���Lt�I���H	���ŗ�t�,��1G�0��h\g(�<P��M�[h�m��\ln�
�3攔����[|�Q�N��ȃQ0�
Ӫ;���Qa�2ņ`��P&_Ь�3'�x�g�T�]�+��j�a�Պ���
:�R��j���*�S�oڐ@�B����~i��F��4h$�E�����irZ�&[�>!�w��/�1���$���>!�-F��ș�\$_�3tlqbl��"nGFcY���A����-�ݗ��b��<�Z��������/%��O�ޜ��K���&gA['P���ј�O|0]M�$ؔ��"=�V�|�Q�o�ؚ��/�'A!6���6�/��i�d�z�A������3F�3�K5�<�/H���y��)�qe��h�$�x�!h��M=-��	�*���3�
:3�0��f�O�������p���ǔ&����}<A�Ć]��Tq�z��q ���@E��9��c��*՜�-���Q�Z�9����uYjO��	Q��)�ۗᘨ�=ewo�?c��jN?¸.o��C�{;=MP*	�n�?��i�V���O���2z�O[S8A�295lI���Z?�,�1∁`IƖr&�f}�y�� �M���_�.uﴈ�=�4�:�˱W!W.,Mgx��z������"�tGA��K@~���@̟�P�?䘏��Fo7�O��&�nM�^���B�k���T��%H�� ������a��oR/�j��܉��G �n�+Y$�g��r���U`��-o=��C���%{�Lf�k _�Ov�q���%{f(6Ї�ꗫ��@@�"������e��R�K�sr�$d7 ��rVFI�������Q���tlZ*��fC��:2�#F��� 9��
d��޼�����Q~��^ju��[)�b��y���{̓[�Ŵ�S��c?��h�?�ef�t��Ng�4�t6D�����`�@�3\��f��.�D��	<}J�?N�S�Uv_L�!�;��j����5�8)@�0��&ZX�*�C��~�.�o�a�xH�$�	?��@F��pSv�r�Ɇ�\E��F+(��}2� 7V��u��,:�Y�O�9��������e�w�Xn�S�t���cF�U#�a��d?�|V��7�p���9��.��k4��/�j����D����qW���QS~�l'��G������/`Q�AB���^&Av��4�Y �3�$l�C�Y�/�á��>�����5�k��1���v7-�x���:K� z��E�do#s� ,���-�!*�����A�mT2h��؁��]ʏz/0�s���ϱ=3�bK�d� �g:�4�����[.����n�9�_0��@4o��MCp��gb�)���_�]Į�igc�W�t\��b*&*�+��i>��g'�
��F?�����B��֨UW�qjm��WU��w����TZ��t
�A�a�.�E�3-���c��LmT�gH?vT%B�� sަ?�g�Ү��50e��|�}�;� g	���YBno�)��fRBf�hI��:�Kٛ�$>���F�Փ��XփՓ\a��s�})g5\F�N~��7�[�KUV�f�b6
�	���,��ކp�P�(�����G/���\ڰ���.�5�n��>V����}L
~��&M�A������ˎF	�D���if6�����	MK�R̱6��/W$�@���ՠr��|��GT���(���ń!��Xy��p,��L+J��.�ԅ#����}ZAR��7�:��� K��:�sO�ǫ�MV����)����,�*�	�T����݂AXe�9O7��h�4��cskV�@3�ID�*Z�9L�z�ʑ����u)����~R��o���X`�,}�r1�D&��%1�B��'�_ǌ����M��(��?�ZP��Γ��6=���N^��I����,�9��l0�>���˘,_(�Lv��7散��l��1eF�ݫ5
%ḷ�W<���Ѳ�0���[9����Ƅ������t��j(fq�-� ��_.���y�DɃ@j��,��P����U�Q�����9������r�g��|��
�VY���t1�f�;�]���OK�y�D��)*�/R�S�Ż�$$���; S�W��C��RM~o�\QSh�᧧���{�oG
�P%x��B]��Qq��aKc	�컨lP���JE�w_�6OÄ,�`��B=CL1�N���e���X�_,J�����e�\�բ���kL<�u�hLv&ɬQJ����a;y4e��&{Ӕ��/_�pd�br������RH!�S::��E���Ä����y��O����oWy�u.#�$+��ڲg3�f���Ͻ���?Sp4F^�z[J��c�]_+���ǜ�K����ٟp{Es��/�٬U{u��HהES�#��*�,��� ���=�!�O���Y�U�M���
�RԸhpȠ�m0 �"�����jp�un+��{?$\�����+Ҭ��f��ln�X�����Zz�2�+���9#�Km�]77��-���۸.��5Al����n��:O�2nwu8�a��� Ԗ	keD��3�����h�&��E����@�mM����v��k�x�Ff�0<\�#���ˮ4K�T-��A�~7!;[����E�q�k��SBq�[��/�Or�)��l���??�.#`˽<�;h��
� N��UIy���|��To)�b���H���n���pCs�<:#���*�m�Kv��q�%B�u�YM\}�ք�
��A��9���4�q}uW�����HJ�ׅ�]��~���)m�dC�����HYmɹ/La�?�9�o�*�B��}&_C��]����c����
�t�G����}y_�h���=��yK^u�T�N����#Q��z"���E��*�\6I���O�Ny�N�ω"r>�0��1��^
�Q��J���|�Y(�!�<q��=ZgL�ӿ9��sWg�r�\&�g��_��`ggX�G��I�{���* ��#~U�*�/&p�@�m�{��U���J�+A5��!�� �3{R5���_���QC�]��� �ph�Q-"�N��m������O�x�A�ʢ�68��#0�3#�KR�k	�i�!w�,�CRo�h��O��Z��D���;y���D�7��7��ݿ*�I��]br/��4��mj������Ui�sO��c�*xu�hYn��� �5��0g5��$�zÒ�9�X�~��=r2��,���LR�2gk�
�����N�^�'Ɏ��Cu��� L���A��y
v�7���ڗ`�=���Юa��xp�g� ��CSEL�K(!I�ɭ�`��MQl�%�Ȃ�-BZ����>�����o�W�'Ow䋕,d�Fu�5'��l��b2�]�u�Y�P˲��q��A����.�����x�g!+�e�J{��<}p��vW�*�å��	i(��?�Ķ�(��/�Ej`����V,O8�S@L���;y����7����-A�h.��!�r�|��si������-.DC2�f5�`�6��Uw��yG����:#��z�O�	H�T��-��\"Ü竝�w��G(�e�8ik��w5�޷��o�Z�����	'��B�0)�����y�t})���j��M�]�<*P�.�iL�*jN�+�`�20�a*8�[���8�}QTX\���9�X�����Md=�	���RռSW���O�V
`�����u1���CtN���d;Q��wD��6J�k:���&$��a ��{҉�@���-s��T�{�>iK�ᱻ%mg�tUз��3P�n��cQ2Ux�I�E���̐B��g�W�B������	1�%��JGʉ��!_g/�ĜUV��DD{����2H8+�݉��<9�m�^�tvg�[���L3��p4�آ��F��p�W@'D=��|��X��n~��ʂ��^T$�^�1�_���Ś�vN�ܚI��'����������E�Y�G�V���0��.O�_�^P�F`$�o�7+���Gk��P�$bb��ݳ�4�nM�U�#=}�tn̈́����Z^�ҝ��mr�M��r���u>���Z��^���na��͘0uP�i['�_޻�+L�����"��A�/�u��	�Y�;����r�%^���u������>:d��hz�U|�� ����}�8��JFԷ�~�l�X15]�M����ōc8�>g�UǞ���ZF����L�T$l��G̟O�0��9�gk�9ۆ��%�h,u��5��ć���m&K ���B|�n�U{�b�c�E��{Z:G���Q�7TZ;_���[��AQ���Z!�)��T�X����}<lRWd�íX�P���׸��&�rtbxo�ȓp�m��$F��G:|#l�֮~�8-W��ô$J0ao<#��@J�l-����2:���R�8=S� ������C>�����{
`	�8L ����0����������c�%O���q~r��R�l�W&J�������,��7�8ȿƩ�60��\�cD��ǒ�����^�֚�'G%a��l���E�(}=cr�ؖ����J��|�������}�H+�l����U��=���<P4�������n<�s�%grѿ�L�4="��چ��e�	�v� 5��(fZ��Ԣ[�b>�c��4�Kߵ����,�8Ii�q��>��AE"`����K�lb��BA����m*�x7�=�!�����ܬ��*:3 /�r�u�7�6���fYX�X@��P"g�fꏬE4!���,�l�˪n�a���/~|-j��6��d�3�_a��(�SD��Ǆ��f�-k��I�<������7��>�E�$�{�>}�(����P��<I�W�����U���M����T6�Mh����=[J��U��߶	���_7hm�s��~fN�6mU(�ݐ4�?Q8�`G�C69�Nu�En����B��1���cWI.e Z'6�P�����5��GL'�;Q��+0�+�f��S\l�_���z(~"#�n��`�U<D��ۙ����!�^6>�X�'	�	h���A�Ci�,f6,��>��*�_������� �j�Sm�1�Nv�sw���c�sf5���^�%�/�Z�9U5�IT�`���{��e��k:e1�N�������#nE�qI3��)&��|6�>�5�B�~���gd�MeߞB��^iO�
��I��	�´C�ڬ8g�of,?%���k��@�3T���X%������7�g�d�2�F�,ma����x����&�U��Յ��/��˙��C۷C�&<?��"CP�l����*�#TTuM��4�%��Td�����m�_'XU�?�K�)�c|ñȂ��v&�<��:te���G�C=Ё�YU� �"��5qb�2(`����h��mߍd��m<A���ב�D���L�N4�����> i��Wg�"��E�����*��#�ؽn�ڝ�Nd&��>����{�9vK&�:\8O
x�_[�/.�����21�h�"��0f�\���7g����~���,k��e|1 =~Fe���`Ҡ;�P^�fX �ؾ2l9]��Ny�12�_z�����4�����{߿\��xE�"?K� ]3?7��$������5���[9�d^~DLF{�~�����:>��L)cp���E�v���;U1)��ci����K�~� D�zSGI@��h
/�؍��"P��VuHՉ[lٲ��ߧWP�Jک,�K�1+O1��Խ��LM�E��S|��W�-�ñ��3����a�=V���,w���[H���5@	�)]��	k�A�zE�_�6�.%��us32$�	:=��i�ib٘��f�kZ�����ų�V�c��v�^�W�lO/�6]RS�_��R�b����<��_uB�� �0\C�m���~�����]:����󌮊NR��������Ø�3�k�6�7���zc������j���~m'��yFvՒ�n���9��Ɵ�v��?q�+���p�/!9o0��4�3�ح��'G>�m��`��)���Pͻ�Q�rA�Tz��^aLS��t���CY$��;	bl~-��D��1y]���(
�5�J�Gգ�K�uj�Y@J�旻��-�e����t���e��ݬ�휿��KUa&F6��d���$!xo�md�o�%�UZ�:B���0��V{Kv��/���b��!a�&��]������@ڿj)qX ���6�[��v�$d���e��U��G.�GF"	����%�]�Ypd ���t܊uƲ�!�����d����V�|���7�}���d֥�����4D�LY�ɉovz�+ϖ=V�Yh�C�?|If��R����b,��W�qې�O��e�s��~z�Eta��@�r��#���kd���)BAٲX-!��?�#Ɩ�z��TxI5�����G���v�Ϭ�c�u���o�.@��y���<c�q��5��ǧ�($�DP�%[b��2u�'Q]�4�'��B��=K�f.��ș��wݺǭW�[���"�\C�
H�	����ތF��Ng<��+�R�)���]�kۉ���.7��dM4�F�g)c��� �KϠ��=��*@A%�dV!	���N�$U���YRof�	#1ݬ���� ��=�`1��e�����/�⹍�^Dk�תП���?�Fc]g$M5s��}�b�s;>]BGYr��ґc�"�$�8U܃�N�E~w.M���LLX�°ʔ�n����0�����}� ��}$����Ԏ1$�e���ȓ�-e;�vyD����^	*׽�K�E��F���n�x	��_��,P/52����}-:��]�6q��:��&_��ӂD2�*���<�g���YEbZ̊�9y����l���#�h����x�7�]F�A���J}y��!.���n]�l��c>�"�����vs�x`:��� m����&X������('��J��ʢ�_�'��l>�ܞ��?�)'qy`s���Q+A�E��#�"U?3����wH��!	�ҩ{��'���%0O�+��RO� �\t��%������^���F�g��n�o�M��ׄY�@I��������K/�醭��×�o��t�E2����S���,�����]�'L
e��Q�n�����U����y����9��p��U���*aE��������1 #	_�5��w>a�0����	�F���ǀõמ��ۏe���fn�]�n20h���H�+���+")���mʟ���� �/�:�eh�̲5�%��QX>Ad���B��.��u)�]�]�0��	g]�tv:w(79��Y
��Ϭ�6$1arH3Ad���V��!F�
S��T�G��,�-�K��k�=O�����e��F2h݁5�+�y)@�umo������ɸ)�LȨ�_���v���1�]���]��ȃ�D�<2�����`>��z;%��׬W�[\��b�Tߐf���b����[-�|�J��)�*y�=�]�����*K��ff"a_h�o^dN�c*�8��^
Lck"*p��A���u��X��?u�=~�y,�i�;�ȍ��m��b��~RLI�Y��xZ���+����ߵ~d��.^{�׭��p�e�}9���.�z���ǁ���O�i7;��WB}𫻠��'��g;	�~���QB~3ϫck�{A6��WS��K3��u�PN���G4�$k��[<f:�Ǭ���>�T �l���*�+�w����᱊�F�4�=��я ���H���ܯx�k��*�=�?u���zJ���������CL���uX�.�C��[<]Trb�s8�ߏG����2���ߥ���~F3w�a1Gde�=��I�:$S�����u�!t��L���+?��8��
�g{<�C�p��}H���� ��¦�����ڨ^R�Ys�(�?����mV:�y��fw��[��,�[<r�iVb� ,����H��
�.[]6�Vꧩj�z!g@q�i[-7|�;��_��D�R,pf��7&�w��h;������j�?��\}��F�_7�	ě6��!'#��U'�6�2\Sv�BG���������� ���
��fq�<6�@�
ۂݻ�������CՔ�Ǝ�y?���,�(�M'ܑ���ąXϭK`�N�{�T��-Aj�����g�h����	g��g�2�K�V!�VlO��s�FU6��]�χ�����'.�)Dt(L&�)���v�`��a&�5א�� ���)K�v��s�S���⏗s�����h*�rJ�tCm���r?sP*R��<��oI�F¹g�̔��Fe{Jn��C�H�q�v��[���E%>��Z�����R�H��b߄N%��WwǱӰt�dʕ���\��������.�p���&����a!J��0&�ظ�?��D�2�O�-}�
�[�V�R%�v<!��~�T��x2?�K0o������|�38�);(���A�(����}�<��A�DM
�5_�ׄ�D�_Yj��U�k�Gx�\J������զ�s��	�������G��GuRx��q�$<�G�J,+VWV�SL0��B���o�����J��%������eXoP��q[8����-��f��+�w�b��*��ڛ�ٟՀ�
/B͡�ɛ��h��Z#/U'���c�W���
�;���yz��K=���M�M��K����	L�D���p�!�F��`s�xS�ܗ-;�-*��ϲ:fY�~m6�0.�S�=R�X��MNV�e��i��SP���0t2N�7
���A+ǚ~n�Ր��E���1�b�O��kh%s��P]:1a��vc�S[�ܪ����UI|�G���X4����ŏ?���M�sFC�4y�w�9iY���z!*K�[�<��o&��Ѷh+�e#�9K��� P�SY�b# Q
���^lG��N�"6x��|��gF2�F�`���p}�0
���w��0���_��2�|ߌ�hu�����daAS�G(����������;��	I:��.�{nYJ5�F�Su(Q���@B d]�x�ӏ��ů;Qv�{�)Gꃃ�]�쎈�f�X�:�JK�\�6HG(G��N>/������O����{�E�C�=bWK��%�����9��>p� �F�o6"��+T 	��L��T��^3mąeפ��)���yE�ψ�����҆��YN�#e��9�D�:ΫO��S���t�be��Th��!�@E�� �j���6+ZRŭ�/��4@O#�x����H�� �N�6��7n�(ߋ2�s�֥R
b��F��U~`�snN�'	QR���N���æy|c�G�C*].���Z�2���%�2�9��i:��J���^:?�AOniu�N�H��ld�d�NS�ʢ�O��������-��v�DښC��:4�#1{�ѥ�b���d_�|����a�� D��i�]�������@8�O�Il;'sz�| �^�'�_?�(�qف��'F�&���Z�M+��=S"B~���k�0.�{�C��CP&K%+G[��gF��=�|2�����5���7Vg���p���i�s���%�NjFy�aQ����sHqT�;F�G�R���n�����)�$zߧ���cv)��r�Wf�N��������)�����*A��&���+�������u��Y������GT+,��Оxjӱ]%#�h����ǢPiN���Vin�璵N\���.��5��O׏&�+��ym����U�����>r��"�:�Ԙ8�O򉯑H���,Nj���H�A����C����%S`�j�[B!���l�e���	��N�O��=nP~S!'���2������\�nIjvJM� o��R߭�$C��3�)���iFaG�bz4��0�����b�b"���TV��������Y�YH�T���5<�X^cick@1��ӳ�?�M;	t�s鍍5�]A���Ճ��m��f��"�|���I�-,�X�9����om2bRS)W��e3��k�)U���=���9��������N���	(d��1��(�"��P����), V����5�7Zp���l{_����1��P6�Du�?���x	���Gd�&�2���R��'}�g/��4ؒ4�y-�*|Y��C�����B�^rN|�t��!�|�e7N� J�rr��1}玹�<l	J���d��k��A� ߾)��W���yN�x�m�];y����+��
�Ȧ�w@�_�0AsPh�����^"r���	m�u���n�U����K8	КM7Q�W��X�m*���W��0&��g����N!_���L�=x/���ϖc�0Շ��l��;
��#ϼ�d���@H���{K<S���BR���y���!��1=c���9yɺ{=n+������{�o�IK��![J�����?�:�U��R�pM,�����
$���F���Q��o����-����!Ɏ��4�>����'�ݺ���U�{���@��H/J�md[���ך0%{_��DP �ٲ�( �b��;�� ��!$��i���s9�p0ӷ��^� ��m�Q���d�X�����9ا�+*�eWX�g�>o�gp*�4�}
iI�*����%^�T�;y:+�����F�`�T@�����Z{���ʠ}���r��s�����_&H=њ@��3�ϱ1Z�r7Ę��I��c{�@��`��+kd<�/��'��"�0Y���*���5�r�x;k�3�*p�9��ȉ�Np agbp�H����#�3F��"'à�[s��A~�f�f_� �(X4���˵d��	����폄aޅΐ�\T�΍�/K1I�	��P���gaӇUJ���\�"��h�]7�@�@�ںu�K#~�F��;��-zy�v���')C����$`A��1���XtE4�ց�g~�h�V����`5Qh��_�q`o����}��Ui�����5u�w*`O��:P&����YY}p�|\"8��r۔`0�k�yZ'�l9�Y���o6����!IA�#x��h'�`�NB!�&S\r����%s��ܡ��pxȥB��ۭ�}�7��L��	���'�G?)
z��X��0�!��]|�w�� ��=?��zy��=��\��=�S��Eـ��.�l��s��(�:k1���Y�����}�.��fs?�!ɵ����	W�,P�F��(����9��v�7�G�U>�ȩ�S�͋i�f����d5%�+��`�a���ӿS"����Hq�bv�(�%����TUn}����GߊN�;=�q���1���+K\TK�	ә�3Oȕ���1���>�}���%!{ ������?_n%��L�~�|��M�����{t�|Ƶ�s���6-0+�gRk�-o:���k���iT���J���-Ym�7�ʓ��IE�0����2��j��;$z��9(��L-�c����N�����m-/��rA᣽'o�t��x1M�όݴ�C����+�Tp�}��e�8�(�'���$��������5�]ƞ f}��ّaZl��%����,8��-ƨj�>�,�iނ��}f�� �xC���D "\A����;�6���R�͢��ג�,������(>'�]�7��&AS���pXuP�-����:�"k�J�� }. ��rHReӶ��au5%�E���2B�v����6x���2}4Pp�a
Q�}�i�Ex:�,����h��|��A1�T�<��cٲ#�U��)��n�&��?rt�ܔk�㊂5=�D�Q��`�MG`_$RU�JĠ��%�����:%�z�b��0��_�@�ި��kG&��
ٻ�<�eB�Zs���6�jl����0�'�9J���XCZ�{D桍0��$rڤJ�rđ�z�_���
T������i�F�ɺ��2IU3j�/������Λ�.�!�U����LF�~ײ�b����^@���6�R�~�I<k%��R2��r�{ol����a�ѫgd|mϿ3Z���	v��l���L��P��^�dzl�$fA��-� �׷��(��L��r���}�ri��V.�=N���y�����P�����tWUO�`QЖt�"�^֐G%N�,���A9]^�z���j��:�9�&`�#���1�tm�Y�KT��γ&��s�������U'�Ӌ*eg���,UNf!�D1f�/Z�U�âaV��e���"D�
_��;�2� �0������w�W�i��x'|a��L���3�@n$�G֜ҍ��D�B�px^Q3~Zq�����S��_�CĢ
�=��|�^m��׳�ѐM߽2l�c������v@��J�ŦB]#��2�ԩ!52����l���>��gb]�sDf��-�+9m�k�J��Z`b��Y���<�rKLc����N�N�w�5���OYi���U߁��#'Qer�DV��g��*N�
���;�g%�[
��Q&9���R�Ҍ�[�J�e��g�6��ɩ��6��
�nq��HH#>�0��M�e+�����D�3�b��y�mW�:�A�\�	9+m���X��J�]��_�+ �_q�����W/:�+y���x�1 ������~�?��PU�$OW����՘��Z�Uԉ_�f�0B����Ɏc�u��d`>�Q�W��#>��k-��������X׉�3J Vc�C�K��->bS��\K�Z��d9@�N���n�
z��V�?;%}�
�w��!ע���>;e�l]^B�;�p�̘�t�͏)+*J|l5�(�_�+΄��P�R�M��l<�mX�fYx��u����C[�QN�)�M��_x�S�x��� �MKPP@c.��7�rړ����CJ�ިS8!�Ц�~xjn:�h<���q�=�������������~�줧��H��M�D��GqDB��(�*\�s~��ϖVo>Լ
�A��q@r���+Z���R��{j��|��z+Ɯ�ܫ�OT�ā��\�7�t7�����E�Vw �yH������Fh=u��ه�|F�{GFO T�`0t��R(�ߧ�Q�Z��1JX�u���&�F.���r���`h��F^2 ��{���(���l�<�4�����#�_9<�j2����u0�ONw��1�B0Bo�Q���"4n$�������U:f�/��Պ.gCK�]��*��H:W=�[e"���F����~��v���1o$���|�IsU�D�Fr�Ak`%�0� @�m��V��B�Ï�B���t����3�mfC&�lʸ���P�b� #�b�_�R����(۽(����"���T`3�I/�a�M�Ya2H.8���R�2j`ꈎ!y����>k0BQ�\]�eo�U��?-����7m��xP��X�Sj�ğ�:�䣦;a ��2�=bƯ.��rg2N�<��"W�ļ�[�a�ߜ�z�v�� if<�����a�7��#�����j�:Rj�:po][��� ���6U.��ޣ�7�"j�G)A��ҭ�pk*�~L���� G��(I'M��۟Ų��)7�I���M�n�K��5��"�Cݾ�ٷV~*���V��V`��DH��2W~rW�^��Y%��7�w�|	����(���	�NEc@M�wm��g�?^]��B8u�dЉms�g��j�t��[p��se���Or�(uЯ��&�%)Пa��L�84N�~� $e䫤�UmA��7���2J2���x�Km����:�+��r{�5�yG��y'^�� ���P �m�FQq�2����]U��ު$!���ӻ[�?��jgn/�w�d�3�T%-�Q)1�o��y��j��n�z���&���)�x�f�Ն��d�F:��엏�4�������UHH���.[w8(�f�A�2 Ρb��݀��>;d�&�e�2�,iͅf%�K���3&�)��%>F� Q\v�ZnQ�ނj6xF�x���YL���}�J|�`!*��Xh��r�Suך�	ٍ������#�3��Iz�p��cz����,���	U�����*��U_��ZE�mЈH���էG��g�!���L�=�)����{Ҟ$C:�^�y?�|��_HpAE6��E8,\;�;A�̘}Dm�h����q��hb~��P*���lu�ѓ�o���տڞ�QP,"9��'q퇎�j����Ў���	~`~ra����/����<.�pf�>o�塄��R&���%��h��7��ʥ��b���2%�Wzy�mӰ��Of[�Ѽ�+��=�	@�`.��I��aS��3�)�wպ	��nɦ� �m<e&�g�F�2�@��cr�A{�k<�`����W��T����䓆�D�7=��휂M��3O:Q���:nm��+�_xU�~����4��|[\�|]��}�Y��C�Sղt�{�)s
�gJ���M�G�sW㻹���?�4����Z��̳~ۅ��[�{
5��c���qB�)9ln��6��qk҉���>���\o���ŵ�)񤒶�n��g���zlF~2.y���|��ژ�)��h;տ� �6a����<sq\�T)L{�>�:3{f��+8��DʤT�$��n�_�3�P�Vѱ���;�}ϗʥX��K���5�����`|��{�g��=Y���Q�l�(���xp��K�3τ6, �.�:���Y�
-H,>vW��śQ�bB��&��Ǘn��>�㌙��8Zlh�>���5��C!�M�Z> ���������08&�쬰r��`�G�ٽ&���,K�}��b�{ w͌���@>h�W��2��e>�쥞H�L���N���\s�{�#.2r���?����}��&^��UkE����<�y�I�'���ñW~؞p�[���c!ᜫ3F��x*-l�N�	d6Fbu�p��Rk�.oe���'[��>����BX۔�R$n��X�[�>]U��,p�|���S��e���z�ť�F�SsD�u�O3�����Tj�w���YH���ۂ��#�JH��S���Z*$�?�Ah�s+0)�M/����}��NO`ɍ�wMy�E�]�J�g��_�J*�<�=��?h7��y�3���qNK�"�kJ��>�5��6��w,)+��g��pb8�6Y��<Z���wd��g��]H[��զ�?
�(v��G3E��|9�@vK��ڑ�d��J��ʠyH�^N
��'Ұ%.�?���X�g��Ƈ�u˼��3a� �Z�s�HփX�z%��Ș "`�"�Œn���1���R��qs̲����\�?����ă�������w����N������)՟E�z�t5h��iK�����w϶�����C�9nP�)ܓ7��v�n����D>lpc�8��'~M���ki��_<�U�$�*߫�W
��	���F��xL����Y�t�+��pٝ�`=a%dRe
 �c/��c��x�`�P�Y�hVp�r��C3�@�\���}�֋�<[���
��a|T`��@c��lG���Fe|4����V�Z�ʘ�,�ĳ
G�H��v���2��p2c�z=kN�3<{/��)î��+�N���&�ř��U�� [�f��#�ds�`Ѩ��:�"�V���ʨc���7����22�loca��s�*q��
�+E&��E!��f2�(.��U
�^�c\�u�z���R�%Z������W)܀���h���i@��%��^�q/�q�Sq�$G�ȣDeoѕ"{��sT�:�Y�R��}��M�+}�;��ث��-��I���w�������׫�����Z���Gy�zO6G"$�R<8Fb���E�!�=ӡ���N��p3z��
؅�^R�K�
��Q�!a �n�V���B�,�����p&$��<��p\ ��6V��'̑7T�N0-��j� 9SPRpm���f
�N͆�R������P'����z�^��H�>}c޳��e��H��Ï.	��שt�F%T���dkF�n/��
�ءF��<���B���[�zH��F����ƦL:���_ȿ�ک8�����P��5�``x�ΠE��B����=�/�e��.�}f~_�7G�t��������b��^��s� �9*[3V?0 �2h;+��'Ul�=f)�֔�V��]��$5��Xk��u�$����f]&�Ș�&���=i�	Ɗ�$W��먪C���"gxAi7�c�?�6���	��#���J�.@fQ+u%r� 74\	Y}�g���C�``���C�@V�s0�����5�.��%���	�a����2��$�e�lUK�<;C|��>��&�2��5@?��DWX��L��J��5P]$}z��ERXD"��j@��+� �9|��ȭ��<�$�k��L���js'�Z�(�E�kVO*�m��x��6��Q����u�����L^S��7��[N�׵9��ʶ���;\b^��������O�&�ǎ�K����I�Zs��Ȕ��̦�>e�zD���q���R�����&���-�{�G�:�:�]V��Rf�{�K��=V�~Y��v�6ى��!$�k��Ց�����}�w"�.ujd<)I���)x�lS@ݑ&QL�"I�[|tg�O8��9��]����.Ք�Y��=��.?8XR倃����L$���z ����B{�<;�����!�fĎ�����ݼ���Βe��!��>��6�'��/�4�7g,Ѓ�AW�[ߓ�T�,���\�E�[nc9R�]Bu||������������m�i��6@i���,T���*o�v\w��h�r�;��}��0���S�/��4pF`�eG�Mk�]���Vl�;z�f�az�?��!�sr� ���\��@iaGx(:[���t�t�����"��%'	�m+��v���rVz�^^a�9��r�cQF$��Q�h_G݄�V�-�Z��/yaH�b�@�B{񠰤��S�E��A�.Ryu� yJ�̻h�]o�K�Ǯ O_�؄y�����y~�_x����>�;���4��SBa{�e��D2�c�^F���<�Z����z(5���C�3z�W�{k�`7?��A��B,k���� ���h8�׎[m�L�?QL�����fc�:c4��UN+��B7�>J�#�E�7F�~�v������B�z1��H�90��t_.��#����D$�f3,���7m�N�/$+��!��"�0�ڱ����{�ʪ.9r(�^j�`=b�[����h� �>~��J���^�%"%f/V�T�� "�V�0כ�JguN��5��xEh��p�Ж��,A /|������TB�e_��[�JNjc�4���t��3�������Øk�1U��Yy��?�z���U�Ǘ+'���'p<����v��}���?h}\��gS�6���-�(�> ������$�&'	T�ʗ.�[=n���=���b����*����߈��Sa�C�� �,)�`�Ȏ�P�Ϲ[�l�ߵ�n��A�?
�M�!O7��a]�σD������W�3)�(a�l����q�'>���#���1\�Z�6"�/f�-���l�e8w�S������Vx���GC�;P���d֖�>�����=�^O�8�N;����w��HIv:<;���5�\yid�ݠA*h���������;D��}Ucĳ�*�W�ʹ.�[��T�z�8�;RQR��T�?�b�ɫ���y gBwu�x{G�����嵁��2y��g�)��eM�a�[�YDd'�#���gR���wr}�ZR�xV>������j�1��_� �f#.���;ΌE������LO�� �p~�e؂�	L�jgٶ���ʣs�0�
����2JA�-��V)k��i�w�W������-A�:���=��H@�7�z)�iS��9�~��w$x�ϖ(���p`�h[=��&_�"�	���S3R�\0莄]ë��J�����re��R���3�bs�ڬ��ϋ����~��Ȫ�+��v�g�up%[��AB�7��l�	0�j�<�����w�i�7��(Or���z�ޓ]m�:�YB�a��Eg����b���e�'祤G�����x,�D�=�lD,��V�a<ɤ�+PƱ���!	�Q��E�ŏ���b��ݲم�cZG�AS%����ʡ�����_+�2��}�
P�����md��Ӆ�L#	��J�#2Ӗ�}�j�hG`�#�,����2q��
B�D ����b�n�Yzi�>�B/���×(�!�rm� sr��EG܀�jp��i m�i�6F��q?$�����Ѓ��݁3`A1F������
�h�O't��T1���*ӹ�:��D�3A'�v��v3b� ş(�}��l��%K~
^N(7���WkӔ��Աp2����O�ˋ�
�`*���0j/�<�05�dZ�3�؁�6��8���L�Ga�$����q��7��O{q1;��e�����/��z'T%��2�Q�Gf	\w���ۃ
;|ɚ �5�Wa�.^a^�)A�v���M�K��~qlL>y�d�A��p �)��itG�:��\�Ԇ�캖�?��0e���*���L'0���B�S���,�� [N~]|Y��[)�\�(b�����,�d����ؕ٠ q�uh�	[n��W(�G8�]`�����N�4��ďSM���$���q\l��^���0Λ@������p;���_"�$�"�V?B0f�:0?YZܲ�l�ٹ��_oj�A���^7��:@Iuzc`�kb��&ͯOjof����\ˬ�d��	gر��O�7��\2XN�'YQ�����3��b��q� ��kjL,�pxx�A�HA�>��^r�Ƒ%|5����&�q�6|�j�i�d�G�o��>9�&Y^Yp|�-w��W�ZT�q~����`0��Y�`����S�w�p��?&�-�EǪi+���f��5UE��W��t�=3,m�L�#*ʎ��63��+J���>�`p5t�rFѩF�2ƒ
�K\ ���]aN��l�k�Q��^S3�y����E;Ti����[�C���\$"���6
ص�fE3Ȉ��w�;�͸"��q$��D�3%W@��A�ƽ���:�����fޖЦ���U+�w���o�*ȗ7���rΈ��D?�e�n0�]����n�;h�e+/�w*i��!��K��F=ԙL�-��U['��X�׿Ά�����f�	���H:#δ�E��\�!�Vte�*^���9}�ѤDl�ӲSO�.Pu��{k��h�ŘL�mה]�S�)���U
`���m'�@�*�	ow(�@lA��>n#-�z`A�eA��rn���ݦ+uU�Kw�����-�I,&z
X�����V,aR�%�������]�����OEn�ɷIQ��Ep��R���l�����ɐ�d���}f7���.�����i��c���^y���Ķ~��LQ���5o��o�j�x��b�U�CQPzk�������#~�/o>��J��{��U�2hv�7��=�yy	_�0��vh@2������K,���o�(��"���&�.����:~h=n�S<�l�'��ߧ���2D�Fv]��Z������(W���S�
��[D��(4�Q�k���S��~<"T���@����f/�(ѐu(�Z �01��f�ߌ��H�&4=��Ate�ޑ���_p
����!����8�KD����+�ih���&d��d��nT���?g��S�I�+)Q���@I�o���L�RHn�Jh�A`�U���Sֱ�:Ϯ�r8	4���"��FlDT|�)�74�x4Ty E���k�<�1��(���kb��m�A"O��G�8#ف@�>�Rg�Y��|.H�>�mM�k6 le�w �5>!"�-+TA��g��(rΩ���w�*z�㵈�Pc��#�w^�V��0#ݝ�C��-�c��� b��r3yE����7*�~�_ȸUvg�Ԉ���}��j��"��d��>)Y$���
5�dIY����H��|8ק|m�6����-ERn��?N��+��9xݵ��f�!�<	��_��ƾ��o���t�M���7�fwBa�t  J�Mxf�¼ޢWf�cl��@$�ʁ
h�E6���x��-���S`=�N��N���%�N%�z�����zsC^�"NȮzH�9�����mɭK�x�Ӿn�w� ��@��@T�h�~�+#z8�0U��<l?�u�lM����Vh��"���ȥD�@��t�b)��~���-w����[�F���\/"�|б�E皚�D�@��:Q�q��Z�*{�8��p��!0ו���.y8$0e�ˇ_b�
�Z? �TU�p�F�c�7����b?�Uݟ ����s��}�^uġU��+%�N���r"�S��DZf%+R,�o�
~��f�>�j޺�N�7ڀ>��a��5�p��ާ�v��}��5��٧���D*v2v��ù;o�I~f�'�ϓJ�������8���&��+�y^1g�F8x�'�m����(U}�	���\�f�8,�g>�h�L�}������n�{Yh����"���j�6��Uu���������5���`]��]�Bd�4�i�A^��2��/wNlh���|������	��/�YA�ô$��봋��TS{�ҏ��	��S��W�F�����%(Y�ဢV�{`ߎ��jشDݏt�q'�	4 ���o�ը�6�N=��-��^'Y���N��	U����5�I3h�qRa�?�w�,۫�u^�������}�i	!-˸�s��B>u�ܳ)q(�m��m�A�����u\|f��\TY�=�6\�	"��w4Y�)��\�z )�}�6�$Y:1�	��� �)�T�su+ؑ}��z�
,�0]I��!dW*HT�`�>�e*��GFϷ�3�>N���a4��PJ�`��<�a�z�u펿6j�H�����k	�j$+��~�TZ����|N��5����3A���: ƎE.�vf�p�)������/��$'ݎ�2��h���U���=��4$�c��Qx��W�xb�!!*��5r@��m�Z�����Y��҂ȑ���:^z��x��5�8k`��,y��xXT���M�P���� �bȦ���#D(�&^p�:4�!�,x}�qU��49���ʠ����t�磞y�W��i��#��.�w:�q�4����(����;WǷ�)1�,Hk?N�u[�	�D直��:"�a(�^:�!(rL��291$��p�Y�y���Y}`���+����T2;w]�y�p�X�#o�����G29�(U��#���ٸ��Z���>���\�_�A�G5-l�}N�1*3�y�ǒ�)�z�_,a��E4���Ɓ��Zv>�a�U�٘la���%� �e�=��	�Ҳ�ͪ�r� �a�����G�NR�16hҠ��* =:�`�dbC��� oaNM*vc~VF�H�B�:텷��}��O�*G7m R��(���g�;K�Ch�R�k�n�ӂ���j��$���Ӗ�^x�~��t5�	k\�O���
Z��6�4���:�����3��>YAJ�r~7V��
��O����J��	��l�4c��n#��V8�&�SC�#C��V*(i ��5!/���w6?N���Iń�K��]c�`~�v��,�!1zX��U�Юh^Hܥ����-w�k}Љ���8��-�T&&|g����ۣ��'��"�h1a�����6�ڊߋ��W�@��ޖt��
��>D/�jB� Ή�5!G���jSs���>��^��^��^���ط�㤃Qx��L����d�*
E�(s��ݯ�<e�B�_��섕����ɣ�,�K��isH_
Z���2.�/j;tɡ����?qd���=�J�$���5\�����*�׋6���k�@W�Y:�x��2)׃�P˧��,j[���~<K�&�Y�D��c��#�#@�%#�1Ƨ�#B�� �򅸊6r�ˆn�|ۈ#�|���wD���*2+�� ck��%đ�7����E��wL
JZ�=Z�X<">�Jci�_�e}j-KH����'Dx� �d/ϑE�t 3�8@��[�7Č�����9������C���Is�H˳��9�e�DG_�yws�ZC��Qh-� ��r7�y������k�:�!xo������k��n�����V��#�R������H�S6�[ώw6[,���c^i��pU��Ī�EMhW�\F�B�5����F�����?�@�9�0�IB#Ÿ�yl���K���ޞ���wх�ma�@�ѱі��F
k�4h9E?����=4
�����3-=��\��8���T�1�鋵�����g�C����G�� �^J�x�!�{!�����e��8���
����3M� ��u�=ԡr��8��R>�6�W`c�A�׼�_�s�p7H��y-	��>���� ����s޿?�>*0� =�〫��2���>�0�� @A{_��F>,�\�¤z���{0�SY�j�$}��@����V��ѫ
�Q�.���%M�C��	�}�!�c}u��[v���d���+�,p�B�ۚ�At|N#�{�,-&��'��ͥw(���t��la��F���h�� H�W<�BadTm�S���R����c�
g�=o6�������&��ZvaN��O[���a/9^���[�
�/�U}y
+�<L �e�DHO|��E݁�2{y��(�	!l� �Ļa`�qT}?�^���i�&�2lK!��1`��s!�ݜ2B��2�Y��ܜO9�A��p!��QЏO����v荌��)�<�(��wiQ�Ї[C�It��r/�<L�$h#�8�yϲ��p%`��+�lڃԯ@��HPE[�-����Z"h3�����"�ǽ@�7i*��8A�X7���Q:H�oS�)��UDW]��i� �4�oe򪃐��msy�cbՒ�[�2T���:c&������7�@���f�}JS/�����^���G�� j�Ѹ�Kh!A�{~��k�_��!��w�K����p�S:�g���K�TvkS$8�+9��5��?4�U���/!n�"E��W�4�5�n�nv�.����h�No���� �Rݯ2s��6Kz�'�yn�����2���p}�h�Zs�PY��h��੦�U��
_q��C�i㱿�ZՕ:"�&c&蜃�$<p13�ʛ9$Sm�@*u|��yg�/
ޫ�p��Iuo�Ȕ���=��J�S�l�C�ߖrg <	Rs0[�L4i'�~ot������qm]cw=���7k���B,� �saZ�� ����n�hv��Ⱥ�_�F�/!�Oq��Z+�%p��j���>=�-�>�R��l�jeW�>sp�j��-�yF=����o��ʢ�C���M�wqC���*=q��6��Ɓ�O[6�4�R75t�Ni�'��ǽ�U5�O%Z�D��ٺś���I��ԾM�o�@��g���"�~G辋Dy��<�Hm(���o�G(�[��*�/&�L�pT�϶�Mٕ�}P ��=����(�њ	��Ϟ[��q˷���h�V)��(��<��}*Ca)>��5�βZ�|+6��/����B��ا��Κ����P ��j3�{o>�D̩�`F�:T[��S���E����N^���`t&� ��X�ŋ�����d�-��
Rj��(���t�4��8o��_.��!m��D��ؔ�\�w��^Q9J�=΍{�ʕ�Z�w���	�a{��G>��ig�������Q�{�k�~�� kIm?�&3Biq}��U֡q��z��@t����K�ܦzƫ-�sFG$Nh��.�eˡ�N+#�s㝖��} ��+98����o4�q����&+7�n}�v����R�N�2WP�rSCMv�_7nο]�fy���x��BdІ?�o��%*�vY':�>�K~L�T|k��}Lh,�\���KI�l�V�7qH���,�
߰��r��7O3r��[tihrt���/yR�v��q�vŗh�������:�!S��Я���B���Q-wЙ��Nq_f�̸��Nee>)��1#��,����u�P`U<�*��3���Z<�Pyp}m�����o���韘 ���f'd���Da�zq19�>z�=��ǭ���y��Z�*�8��bF.�MaE�� ���5�J�Rkcԓ�5��Np��x�ѝ0k^6��TY"wTDL��/D��+��RN`��@���L� Ήt߰Tyl@��2k�Cԛ��x�73���2q&S���ɖ���h�޵ɷ䖦��	�0r#Q�����#Dci�e�)���z&�>L#_l�P1�A3Y��P�͂A��][jxw��u�qBSǲ.j風˥Y�E-x�Z�Au��yH����b\u�T7֕j#ȩ[yUъ������D��iA�d:�k�JG��V�Z\��!a�v�n��sK`�m\����[JI{�U��`hM󕛫$\�g i��S.�LQ��B�w	�ټC*���}m]��5 ��g�-E{�p%�ڪ��M%����$t�RN�"ⱴ���'/RX����qi�Y�2�N�`��ҍ�~�#
��$#���d1%\Y��\�����{��p�1$�$v�ًh�?W��d�U:�y���:VհO�i�u��#���EgG4�z�q�d�I��M��+��YY=D���ÂIMW�`,�}��w`�
,�x�޷�K���[>��P��B����qݽ|d�s�p�R2n�}W�8�Y��Y�E(��܊6;�,Dt��H]������qo�&!�uy��e�z;���P
*8��IW��M.����1~BA�L\�%v3H2�0�%%��ƙ���0�D.t������v���^�?3�DW�e[=`��i�C�6�|K�|�e1'Wː���r�ʇ���%Ґ"���K�zR�3p�Ѡ��<�R2XX�!lI7�՞}W*��pq��tzpJ���$_~�H�G��ڹ|�Q��Dk#*�������ë��^��1���/
R��gX��=.c'��b�X��S����TbÒM����	� ��y?�Uf�P����ͼv,OL�G�g���n]QC�@I2w�`O�4��a֭�;:�[ yNϻ���W�M�$�v��c�X�͎�x�mP�\�o-��B�u_h+8�btx9�O�K��t3le��U�s��Q�~"������Фz��+�ߦ2�{��Ru~Sk�P���L�{צ��2�$'_Ʊ!����εM =�o�vGw��2��cz�
��6F:w��R[_aI\�=�I�R+�4�9�v&ٜ�="�-�-�Ը��5�a�>G gm���S�_L��+1 %:}��aO�2�kx��ZSC��\���2�`E�S��1�,�r�SI��!_� ��L���w�RW��v{ۏ�n��΋K��*��	yl���r�w�i�m������]&Z�B6�����;��H��4Dn�Q���	XL�#~�Aߗ����z�zɋ%�.$]�}�n�>2��# ��G�zW>=�i㐦9MĎ��$"�WZ�M\��(��xoUc5%D�Ƅ�˰V���|�n�;B
�A/�W���Ԏ�X��f��M�7��/���:��f	�v�ؖ�������y�z;l+���VO�ȮA���xCL+�0;�t�˄ГE/�Fw����S���b�Wu��C��$���3N �H��J���N�f�h�YwY����醬]"y��D�}��q�7g2
x!��rzM�0����ɭ���C��M��n�S�gH����XXϓ���a��RZ�T��B��b\����nG���Y]N�.Ìi�n���O���)Ȅ�B���H�2N�IK[�YR��'�:2'Q�P9�{���jp�L�t�͗�pxR���0�얬 ���b���O������߸�0�Ӯ�1Y^��%�����rQ]y�4@��Q���[�d��}���(a��J�d���;��O�*bY8���B�/���k��s�f�.�M�hBb�|�)�v����Y.a�KQ��{�Ro���5-��f*[�<�[ԓ��1�ԹE�+�ѓ���ߒ]n;�_�c�jj�M�������� �8���Q_vO�ɦ�@oU���ZS��?A�.�Ə�A�N���/�(�=3�ݗ<�č��-�T�B���S�M�� q��զ��9i�вe=ɻ�xP$��@���<�T���̗KX��<�,���宐{#�%�\2ͫ]�����Q0�x��u���2���s��k�J�9��UTf�H0�S{����Y ˟�i�1O�8P���rĴ�u�߾�O�j�� �(*�:�q��3E�ܚ�� ��w|��i��04��>k��k��>e֢T�VG���~��U�w{#�W��H���ܤ���	����JAʳvMz;�f�%
�s��~��`��γz� �q'*�a�,@�pռ�"܈"~�t��
T�����Bb^�m��=��jq�x�h��a:�NYսQ�d�|��2���߁������ȏ��G �D��j�u�r- �����ܯ��=����7�ť���&�v�����3�萷d:@�f	l1���w+���hS8��y��}�Q��d��
�+~42[[�p�\�s��,J��2X�kR��,]�ͅ�N7w�^D��~�D�����p\8{G:F� Hj!�_�o��I��N��� �Xν�J���(�#�ڤ+r�֒d��-7b9� �P��~��?p�,X�1���v�Ї��%?��څ�еML�W���=���<�`I�''5,-��O�M�����H�qN����
A@Iu��u0����M�IsF�6R�	XN<���C�n�	Q{'��GOXB�A��=�E�i�q�e�k?#/0N��Yџ�vf�<f����_���NV|>X�%TK���⳰ ݣ-op�����`�w������K0�a��*�xψg�F�r�%�#�(rL�
6��V��?L�mh/�h�l�5X|���H����LL.�=r��5��Č���Ƴ�2�m�C��4K �U��\Ri�ۛ����Ǟ�A�̨��(˿��b	&;�Z�w�5)͜t��9�?ۏ/r�v���CA���
<NA��NF�KVKsj�$�/'��o�\Բ�����Vv�,q��d�5%#��61�c#���Fd%�%�AE���I�X�ƶD$���a�G��"[Z����V�I��i٢��*�O�u�8�2�˯((u�W��JM�fgͧk��i��#,��!Pl�9f�R��8~_���BJ�?d���ؿ&@uE�'9�2>{�%F)�E��e��lc��*���y;���ʥ��	%�p�%CJ���N�,�yD:6���5���LL<�3$�E��f�����V���'�{���<30�Oْw������(�ޚ
'�M�f=+���;�&.��� 2���J�!:���#j���1�8�\��V�G1v�32,���J�R�>��O����q(�ˈ�N�����r�/ck���j:~�bΌ���p$'�z����KV>�/IT���'���m²5H��g#Ӿ�LB�gI����*�RF/�lK�=V�%��J���Jȅ��+�yvy����DCqC��F��_+���ô��@R�|�� 1ֹq�]}�!c����>�,W���岶<��qy����z�?���� �R��X[��N�"��cA�J���^�M�ʇ�r��Ҿ��yZ\�ڭ~�!cf�.����uH4��c��g��&&���SL��Ϟ�>���CF��5���#/ĭ$E���⓪oN�X��h�x���5�֏
�����Ă{��o,�r�S�\�vy=���=����I�1��~s�{��!����`�5����I$i-��yF�����>|7���@����2В�T��,��݈��A�-T���	AOO�^aeܻM�4�6���˒��/%ߪ�8�4�u��F�4��1��ju�|�=U�LPZ)�s��~jo{E��)ƾ� �wh"�_�9I�|^O�4!������ b��xy�P���3�<�;��}��}9~��l8���A/z�nc��Q�?~	�w�T���>z|�� JO�ݑ@�2}��U|��'�wv� ��6�[�
w�#���;����t�~��QE���62��W��G��{+������N^^�o! �u���.|R{( `=r���� V�Ϛ�d��d@��2�gǧ��������hd�_��sƷA�X�Z�����mK�U�/p�K�:-��8��.h�!�>���y%
��<Gon\����9�Z��me��j�{0o�/�zã�'e��8�VBB�S�6WX}�0��K��l�a(�����sZ���8O�3&aq#+)�X3M������g�z�ׇ�؆=�,*A#Oz��WY�K��E�]�ͶC�<X�buv��46kޕ�:P'>�1��QŇtX�{�GuE��㴌b~G
$���LF&�z��?�Mo���(�:�6|� �,�d��O��Bl�"�O�j�"G��*�w�X�����k\�8
|T�`��9QMs	/[�{X��XΥg�MB����D$���FFG/n�%c�a�S>UD��G�������$�9�ep	�� ���p@���ÄԹ�:AE�S�k�79����y�������{�&��[D�:>��#�+瘗�X���Q��1�i����#.�s�(��Yt���6!���+� ��5�^���-O��-��{�W3FK"��OA��#�ӛb����eЖu�;�1���D�
G�	�PQZ6 i	��úa��(lZ=�
3.<e��G?SK��D�.+"�bǮ8�$7�׋:Y���ĩt�!�D�8tAt�K�4���X�ccd���ۅ������Nh\.~_8� 7D>Q��C��x�n���F�c����*�'��m�VWϜ���#����y 2�O���=��5��j|#�mR�Bе+0��r�i�Нx���S��̀)m���*�e+]���<}�q3��>�:_��[-�V�%z���_�N���y�G��l�����C�/4,PZA]0E���`[��~v��v�r�� �˙]�F�CjK����N��A�p�p;pӻ�Sc������T."������������]�:�ŉO�&�a���d"�#R��V nي�E��������LsSZ�x�����\)z����D��7�������_Hc��<�2��X�G�y�{��?�.CS��V��$�rl��p�����'?-��Ay%h�vP��=K�4O<.��z`&)�49P�LJ��&���hkZ�x�a�+���c�:WJy�g@�2��4�8�"�'���?A<���w}k��g��8�L�z15���w���̘x�`�ZF���&Kw5�<��F��S�Xvd��wuw�=�>�G�c��C=�4��]Ch�� Z��ύ$�#����@������i�\��Qg4r�y������'�������HcMi�G��'��w�jc�慢�ji��fk��WA3�����/%Mi����/��=T��HQ�?'�CGl�i�ήf�Ԑ��%�[h��v��pj&[�-���y%(���Jb�r�#�,����{��U��z9�����}7=?f�J`�y��r%R��keW��X�τ��/�˲�,)=��p(��P�3	 ��z8!��x� �.'���l
 ;�ú"9e��ZRzv��E���� ��$sg��BS7�ff��ݳA��c�@qI�Ox����0�)�/y'����ǘ,��3��i6�j��S���S9�`G�����_�� ��� |@w�V��ۇA!�<�T�+�1�G���(�ŵ��3���~�����{�Z,���Zs�h'o?�O�\��^$����,S�qH�mX:�ix��C}t1�_�_�������a �I��e��z@:t������;��}��D	���G�2��Mӄ��˱8@J_$�O?�X T4,�C3pK֭�}
AUCj2\�(q��Ng#^s��Vv��̈́s[wc�;f��c_d����� 7�[��>Q|]?ұ�T� >o���,�;���%�ԟͫ좴�K4@#�+��Q��g��@!�Oleo������X�`������5%�ᤡ��"�GmR|k$���|e�t��=nk�( ��|Z�쉹�FT��@!��.W2�rfx$hN.U�
�_G�G�Q�Y��2�|�]n��Բ'���G������?(���37Qʌ�w	��9�/���2%/K������3�;JfYY����$ ��8��ų�?U�q�	�31�v��m�j������A��[Vwh�?�kK��]�xix��S+�ڥ�0� ��L�뿯�O�0ߏ�W�7�NYwB��ٚ��17QapQ����ޑ�_ƄN�--$������ުvH�q����b��?s�~��;�G�yY���}������O)�w�4�ȧ;6��F�:�D5�ۺ�j�oH�Ib��>�գ�@�j�9�[�w=��u��=�'����T� d�80J��~�1p*~�*����T�Ч��`��ed�y�o6���}�*��V���Ӷ��fΙ%_�vs��(�8�]�M2ƛʇ��@����NF10�p�l��3�φ��, %c5��F8a))Ԁ��D�pE���e0IJ~0M���~�@�O��� aց�N�_(O�Oq��^R����"')�ʃ������N��p/]��i��,�~�sP#�?b+�i�2AƁ	&��QU��읭B�(�z{I=)��z���Gt���V�����M��6������rv��Tè ;�|�p�]��B"�Pi��}}YeO�Cm�\ ����Q0l��ɪ~���,�	�����:�v�'�#D� �����<�o���E�oz�K��b�|Le��.w��� P��#��Hl��v01�b�&�˥&B��*�Ǜ�'3bJ/j$�)Nsv�p�smѨ���-�]���n�@;�H^��R}��-֕D��3�D2ч����[tN>;,�u�OSAH��k1׸��`j5t�Ga3���P��	����_q�Wc�X���l�/�JF���
y���K��*���!	U)܎��R.J?4���]j�*�$.&븗mM�C|?�}|{wV�']�m�k/6�-}/�c�D��
UY����Y�޲�SN�u[��n�����u����{�L�e�ZDW�G%ɺ��� ��T�ŋ� }{�&?��Ȧt��q�+�������s(Z�Ѧm�N�d�ZlF�{���I�E��>�"������]��:�z�趐�mگ���TT/F$c�ɲA@6��$�D�����S���6�ƛ9@tΪ9��Nɦ��8
�E+Ƽ��bFn��r�-7���/�ˠnV��,���5����13e�m��L���ڲZ3�iE������I��VS;��4%�7�աMu�����a4��z��{�/4f�;߫�4��I�t��dT�\�i;����ۻNH��SC�9F��y%ުQ���c�..�0���a�°o���ȱ�Vr�R�}���r�L��Q��2_ո��i��a���a���81�_��21`/o��3��Lc���h��^(|��	�|����C7��y���$e4[w�N��W�jh����*Zz��\""k�[�ΰ'u�4��"&�T����w��w��]UdR�i��\x�3MAB۰
�M���C�~\r6J��IBw_e��p��3����'L@N���<�[�����:O(�:��>k�c(&����Yٲ�-[Ԯ(%2��Ǐ9H��m�"�&͵�w� 2B%�$�$��ܱ���b�w��Xf�(ժ.�Nr�1-��Zk'����̥+Ύ6>�%-~=�'�^c��d��bRڦBؤ�9JV�)Ȍ5i�@`g�9��;FO��������y�_!�}? ~��G,6lA���ii&�у �����4�ꞛ����Ol莤�d����[��|�HŬjP�(a�K���GD��Q*Ǹ���_���tDvj�*-��]�FPr
ݣ����<,�Yds%vJ`��̻�N��,&�U�(���YJ�A��H�+��k(��A0��4om��#%������e�����S
����5��@����$D!�!3��U��HV���(1OL�NBf������.T�H��~Q���I�7�]�FQX,;/��;7�N�Q7��.��uT,�P�R�7vɿ��yJo�cpzf.?	�e����3|ۼ+Z��v<�LF���m{pq����d���6���W�>�@��o���OS������4��sp��ա���-�9�9�R�RM>���s�WH���^�	���n_�9n����AU��ǰuJ�
�ޓ�^d'�'��˦/�c#]q������և�t�A����z#�x�1����c��2+z)n~j6-���mM̏������*r?Ўl|���;#���fY�-�SNF���Y٩Ի=S|y��"�Y1e�H�T��x���9��,/����"+B�m�:�g�����%�d�X5Civ�=�OІ�H�X=����v�L���^-��y��cĔ��G>�k0���I0^��{q9}�9���5��e��	�
���i�?�2�^��x��(ō���p���5���{���QM�$�Ή3;�9���a1�Ê�=��6
	\�l0�~_����:�ڑ�.aA����q"�8��y�M|6�(��se��i%B�AG7�w���:D+*Ĳ�k���tA��A�[���gYk:�W��o�8�E�O��(�`��*�]IK��e5��4,Ԏ�ce�2�6����e�����'�:�q(���|z�+�_��:���ԗ����ۏN���n�-$�J#���~�@N/�dܥ�r�f7������pg��X�#
��z���O;�7<�27����;B��\
S6���V����F� ��>��3�{�Fװ�Lf�Px`ʷ�(.�����c���C����S<\&��4w@6��kʳ��HOR����4DWd�̌�� �U~ݭ�p.�Æ�\�x�*4m'E(&�n"gZc �d���jH�s���1UA�a�Q�8��*r�!�����R�-)1�{�c.�/L�'9�Q>r�ƍA�tN�C�ZR�p~;66�ͬ���; �=8�<��-�
�.�α����,��B�8`�&��:=+��I�,삅�-(�w�}��Lϰ����&���աx)͗�����o�5����j�/G��Gӣ}?Q���T0C���lZ�Y}	��z�Fr�*���ldTXi$���J>iF�C(\婎׊�f�l@U��,���\IN�B���[���U�l]�MĪ_�@�f�ҧ�Bw�!Z����|�-L�v�A
�v:U�^ ��~Pج~�]��HT�T0wε��Ԃ�"��9[l��@r���Q.k��_V��&啤�T՚�U;���<��N��7�LI��l8s�=�����_�Qe��L�F�z�,��%���Q�l�N�9�Ҕ�N��X��E�`$Am���0�j���5�Gv���W"E(d|�<̓W�h�8\�3.V�5�pCҪ��\kk�l!jv�q�c�iv���~�n΋�{�<5��P��n+���􏶂���X}/yS�p�cu�8�	w�l�˾�����jJh���dQ����=�!t��<iMy����@��,��MK��к��g7t��7�K��!�]J&^~_�M~��ȍ ��(��^5v�~[�ɾ�px[����6�T;�5�nk�%}���D6�u+����N�����zk4���D��I�iY71!���r��W��$�CY��B�`���G���$��r��7���:��s�$aF	���y9�kʵ5d�s5'���	02CV�8C�#=������&��>J-��kK�A?ݑ�[i�f�)"mtM ��jݖ���� #��ϣ@x����e��%X�l�R�L�}#�iGx�n��3�*�#	��:.�!M2k���;�q�Rr�h�ݝ\��\�%k����y���hfJ�+'�2J�t#AO`*��)���B!����YK�ZT�c���_=l�)Lܞ���&S�R� �dK��~�"�َ��D� ��X�LQI����R��?��+4�����
Dx�}rl�/�mvT�f�\D��Y쫝SkX��NBg	؋��;�!ق2L�p eO��AW��j����dIYA�`�_Ҡ��ڡ����:� ���S'�~��w��ӳ�l���){�݁^�>���>G�8U�&��OhX�s�GP�/}�G{�h��S���7̄�-��&��<���a=�7���9͐�=�h���'?W��GG��FNe�����H��A�/��A��A���2��#�#ڔ�͹�4�G\H�{Vs�6j#�w�?�x�����r��bB�-�J��yu�3[C�TRE�U�<��H��޵��~&�|�	R?��������8{�ᱎm�닺�˸�)2"P,٩���ъ�a�H~��rjי�B:�߶w���-,ϔ{���<�N���/��^��g3p���0���#���#k嵿�G������$=3|��EiJyn����?'��XUU���Y�)���=?In�6#*�!�ݘ��,<~��R$-�K��w�j-�|_������ٔ��9&��
<�����~rÌ����|̔�d��6���$d�5���E��5�2�S�G����w���~�Ƚ�+)��i}��v���[���xP���81���|oBR��Z6	7� �R��T�f��-�
���v}ǥ���]�9�ֿs�;J~�F_NK�t/$)�W#���ދ�:П��1q�����`���.�����`��a���Xz�&J�*bKdg�%o�e�Z����O�a,r`�����^g.����v�0!f&�
�����X�u2��������=�'�VWSC����Iݘ�*LQSCdK�#�U6�C��@c���*��iW��� =	�Ұ�����Gj�~�@{'K&Ӗ�D��fK�s7VI��*��1���1�� �0WPB��ЅY�F�&���̸�9W~ �b�P5�/NTU'�����k���1�E$v��ZU�˼��"��J�v����jR{j7�L���:�6�q������g$V����.��ѫZ����cH�M�V8ȪU���E��H�|�m�8l��N>�Q��0�im�a����Ht��l�@?��#5+]`D�Ų�{'e�N�V�u�x�k�`�
m�F������Jmhe�����b�R��g�扔~J3�E>��� �T��Q\��9k�a$�
���@�����zR��d�p����(c���_IHJ��$@��%a,�m�(��4پ���
�L_�v�Z�B�bQ����S�^î�/Ux�[n���A�a��#�D��i��SĔ���I$�5L���au�x�L���'��X����Њ˚�"��{�M��"��t����4	�>.1L���l��=�4�&��PV�Ԯ�j�S00ểq,���v��.�A���M 
��qIy���P�����9Ȯ=���J����J�xGSЗ�x�Z���d�������F-�g�K>{վBBp�#n���p�:��Y��Ill��f^[�[ҽ�甹�PR�7/!C �U� �����kFr�e�`������g��Ka�1�K���VT��*���z��3I�r���*��U���_���/��M�re�/�B��jD��u���F��"!��l?qU[���-[��G8c�e�`@O+pJ��4p
��^g��sEWZ�%�䋢��fя#�><)C: ��;�=��h�p0l�K+��Ql��L�b�d�&/����� z�B�!�:s*yЎ둨h4�ߐa$N��ܡ�l����	sRc*��pWB�m��hH3-;
�MS���j���qo�gQI��|7�#��>�kT��")+��,�Ι�hP��vp2W�	-^4&�Z���: ���
������\����k&O:��V��Sߤ^�H_6�r}v=�s�;[��2T�8��[W���-M=B\�{�Mh�B5B�^]�)_P�����m�o���G|W�,R�d^kzj#,����Rj[�v{*����t�$zW��2J�����G&!'���c16Y���.�����D~����;�����x���m,~4�`�j����O��������G/	�x���V,�����"C�m��	M>�ߎjǌ��]#�e�s�Z�cWYDx���^H�: =KI0��^`l�!��ASG?.�����h�t���� ����AYS(���0H�^�Kd��s�qkے(W2�k�v�,�8g'�آ׾�`�ʶ�<"�9a81ą��XRV� �f�R�M�/Z��d��/Eh^�H&��A!��/p�=;���"B �
K�B>�^ ݀�vѨF�������%j��9��l;=�_�m��V��~�bdl����,���׃c��Đ|�i�sD[��gj�dU�ċ��m�*���B�	���?����	t��z
�`<�4ב���Ň3�=����b�nb'8� Ai��G�� 0'$c��h�Y��3��Q�~�1��Y�B�y���[TS�W<�>��*�����Z�V�p`N��-.v�2�nSLOU9�	g���2����Z4˜~��a�M�]���[B�m�8:Np�i�݉~(���aA$��gi��
����8�����0y���}9�D6U;��,Z�5֘�D�<?�u0,��C2�ܬ󴑙5�T�
�F��p$�񘱠�1�����<�Î�*�"ƹ�3T��y���[:���'�#��3=�\��Q���^��w^���r�ߩ"�3OI7mh�����3+"U�c_�^�n3#�PF��4��a��>�r�y��!� ac���n�oY���	Ƶ�@9L��E�1�F)t���z���4K`���f��M̏yn�6CB�T���/K�k�ڀ.{Ta3����!1�M*t�Z��V/r�@ �ۣ����p�/��d�lܡV�0�#�M��+џ1[⏢=��
�)���>��4_��uC���{�����Q޼�pDq�� wRÞ$kCR(��H���Y��77884`@�7䪫�����+�"��$Vg��^:e�ѥ�h<h��dhP��Uu�NV&<,��`LK�R�LX���R��t���^�?t�,^��D�Le6���Q��GRC>��S���&	:JlG���Y}ͭ��5�&xQ#������B(&�0�K�^�+�n��K%���ݬ^ć�K�N�d+���t4�w=��L�u�		,�L|�&��Τ�����U��-��N�^p::�s{�8.���jۚYQ���S_V<6
�~�}��)���+#����&?e�ۼܫMd?���ahS1���G;A�yc:���������)���e�<9��E�@�K�
�Y�MLρ�TT $z�AI�Z�"8�V��T�kTǶ�b�լs�4�\�ٰ%��>��mA��NMofy�L���X!��F����t�����t��3/8۰[a��
~�ժyE�����ީ0Tֽ`.�e����s8�!g�6ߑf��8؀��E:���_��\��6ۍu�,k�2�V�4v���ׂ����`�c^������#eP�bc9k{bw�d��}��ΰp_��*8�ipҎO�[T�&�p���i����^~z������̎��n"x�#AL��Ì�-����;C�a^��m��v��K(Vg�OĜ�"��V�y��C�5�tS��&ry���2F���G�KD�{�\Qr�lC⭳^P�j77��F(ބ�Z���g@"��@#���!�'�/0�io#3W�yՍ����1���XJie�������7�L�N ��U�5���6�*"%���v�`ډ����$��W���4���X��0�?���&]�<Ϛ�KWSO8g��ŗ5��>�w�F����I+CV���7�z�Rਈ5�.D���PK���{�8���T��mg�+�����'����"�f]խc�N?�;Ra-�>��u���E�,vv�S"F�{�}����^�Z�� ���yh�n��[�ߕ���ux�v}=n;�M6� /�أ�k��I�X�qlF�A=�b��������n^�)W�����dw����˩��*#IkΚ�7�d*Dd z:�W���3S)�g� �'�wą\����@��J�>��ߘ���շC�S�kྒϕ*-kq�'��t�{�<�d��=�!Z���N
�S�؊�������ŋ����W�ݲ:�>�x�1FU�\[:��S�� �Г��8�H_�MLv��X$X��[r�J�3�=�_��+vP!^��C����UP�|���M�^�-��s���7{9��zW�n��A���<y��q�7���5�}3ϙ`ſy����Ɩ�g�ZҲ4|	��El���NA{�4��]~�O^��`����8)�Z�X���$��淚���<ۿ1��^��"���N�ϙA���-LǬRkOD
�� �E��H$HZ���r+��g䣱��� ����W<�HzL[��m;?������6�ݧO��R�W��Ɇ�XZ�_K��X�p'���˯�|NV�;��E�߰��B�����SJ	A��n��Ec6{�\�mG@H[Q�}�j46��L�Lh}c�n �oӥ�@���������g��mѺ��d��D��w��\�����b����k�*��٧�9V�KΟf7���e 5�F$�������`w�$�"��4�:��}l� ݮ�j�؛l^���#,S�����{901�J���X���뒳QKy��#E�[���ϸ��)�Y�sX/�ڤ�P�+wpJ�}�K���nF��ܭߣ��|�|���1�����9�_�������ē�^�+LA���M; Dbm �g�O�y���gn!�7�SZ�c�t��h�_��<4�,�t5��������P����ꆶ�n����
�֔�в���@� �8C��r��+�64���MM�co��=K�C_�xn����2��`�#c��f�L:�F_�� ,�@�>�X�|.O;k�_Z-}nИ�[h�J��C�Lο�hݭ��EE�<�; S &�r�޼�/��X%y_(���ciT��tgUV_6���fr$��da-o 7j�¤WZP�o�d��Vl��1�H3���	�C��]w D��{��w�e�]0��G�d��o�8Z4�{��V#��-�S
�W�*�w���S��������X*�� ��%�� l�6ѵ�&���Xfځ��LX��G'eyE�ga�&��cR{�H����O75��]u�ERP��FCQk�r�I��t���yA� l�J+ε�#�b?v�w��&���08�����̖��ٰq?,�e���)�o}��`��"�=�gm0�wo����
��zr���>�ֳf� �-nBkf���'�������4����xB�{� ���T���#"���v��Y����.�� ��q�>ؘ�����0gTT΍;10"����O�����7K��'��mܳ��/y#�@��2��Vq��ވcF#�nK��zKo�g�`���
���")@% .U������7N�~� ��4;w���
lې�lJ�5o���5#�� ��@�Z����E� �C���i��+��;:�|^���#_�(���"������X#��&h�AV�&�C��[%	.��ۆ����>��?�'�ed9́��b�����I���ωY'������wv�C�r�Th�؛�,��t�-�
D9"�O���~��zγ݃2��ҙ�&�כ��f4h2~��Q�}${�Z�+rbiN�hC��W��8g��/�iK�{ʁ�\����`�"o&y┤�f�'��H.������{��I�㭛���gO�~?��R�-�C����R#d4!O����=�p;~���D�];ms�A4�~���t0�x'w��K]tx-I��6^ ��yb�C��ob����%��
�Ń�T��SY�UM�S�����sDm���~�=�rZ���R	�C>2RQx�h��0��MB����g(�n�Xg\6)���X�[�e�0CJ~�vm>Q�����I,ƿQ�����k�U9�p��,rX��ԴW�K���@�r��b�����(mR��xv!؅50�����7�c1�+&��Z�$N'p*�i�eL����ai�O�ӿ�P.p��0g�!���H#hY�CTq�&��oOJ\hz�D������po����4�o��8���q�q�V�~��ह����t4!;g$	ż7��HPa �1�RM��<x�l���K'a}��QP�M<�u�?}+���,^����ltY�:`m4ة��D��C�w���"��ȥR���͑���V���L�F�h<�.�zڮhadk4nJM�����V��Jm>FX��ţD]]�\_xN~D�a=�TWB��-)Ax���4��Ľ�Y���0�~����s�Ⱦ
c.��!��
�@��p�p���P�y|Q|X�
k�X �];0�J&��W�e�,u�8Ao����/��w�͂<����<���:�|�{�!�����)0�&�c�L����ȹЀ�6�k��~���6��Y����2U�YF����c����|�ペK����C쵀�j����m���p���.#�(u�\Fׂ%��`�sI�਋T�$�g�̖ ����fj��<Y�5�T�M�_
�w?�	bx'j �RBP����KD����y����_]�H���\5�惸����4u_e�[�C�}�O��05��f��2�����"����J::l|]hZ��gղ/�d���{��+CV���6@b����(R��W���gEl2B�@m���#8��J��7�g,��I�&!�QRHё�}`d�P��h�au��t�.;��]ȏ�8��֩<@���X�sg|�{�eW��;�}�q�x(ҹ������UP��,86��	��y� �Ƃ�N�*
�9
@O*�!!-1f�`Y���k��Y�Q����U�j��``\CHz><f�xш�@|P��7�����c�T9�ٸ�i�9�u �{7�������-~�+��W�Bh���8Ɔ?5\����
�FA��IX�j����l	Ž�6�	�T��;�^��M_Z��__�1RIW3��2C;= |E���]�T$�����3	f�e����.�6��+�f@�g�6
�SB�zD�mВH�B���K�9Mk���P��W�\�9�IU@���,p5�a�t#�P��(���ε�[m��6֬{9�S�k�ӻwg�_�ʌ���Y]JY�><�!0��;��h���x�6{���U ʏ)�e6k8��(��)�p`e�, �D�Uyb�_�_2�{Q,L�58����/X��?��y��P)ix��UzԭP���2��+���鼋<Pۊ��;*OO��{p��`�<̤�t�:��[�
�d�ꂌ�C���dA��	1��p9\ӯəC<i�E���5Z�L(ŗ���S��EU��p�
d�=C��G:���bY��m����s^c��ǖ3�32	�VE2O$a7MD��k�gb�N	�H��������������Sv���'�o�R��f?X�̐�z
�"
�G.D�{���۳�?�k���XI}
:�\$�/���M�ڹew�,7�V�L�ן\>NP���I�*2�FB����#�W�[�ga5b7.~���}Vpn���ƜČ��Мr�'-�§-�o#���_���P�TC��G`�����ٯ�)^uׅ�j>H
�<g�������a�~ 學�;1��ب�U��ȭLY|�ڱ�X���fj*�CwB����O3��.�豞���s�5�P�1��m.���"�nI�Q7����P4�γ[��|Cg��pA�6E���1~v<DƦĠ��ؙ����9	A�w5��c)F��E�Z=!"��x��)S��4a��?���5�֓'2���/7�v�1��׿���ŉ,���@:�2cA�i/���LZ�/�԰�3L�x�>�|VF�5ؼ�tG/E�M':�J��f�}�\��>����u�D2:�GԎ���7���p�8.ǘ���
^��¦w;{�Y���P����}�n�]����m\�J��bm6enƾS|���$~G���e��B�.�i~AI��(B8�>>^~J?�p�����q�ẓ�������L�GWW��44��2��D>�K	�fRU��'��]+���A�.�1����K�]���M���$+?Yo��o�Ս4�D;~��t
,�z^�'�����U\'�Vq��/F�B�B�f�����q$�W#��V&�Z��g���R�6�}0f���?P$ޅ{�"릚Ӽ^eF�qgx�Å:<T��f�������X�	`�Q�%��`&߅�l
�vj)"�6B��K�wb�x�Wýɰ$�YRssS�V�F����/�������&��79����>���`�1fVaM-O�K��@�>_~��b���.z|P+��x�)�@π���?ÿ��c�X�V��Q��Y+��Z ���H��ꧠ�
��a����Il)��6���/]��{d��!�V)�\Y/��2r0�NT0�EW�@��q(�e���u��Y�i���9��JǼ4M��O��-8���L�JD�X��Z�bm��neG���̦��tmM� ��*@��،3��2���ؼB�V�dmC�9��h����x�h�`�k���-�b���w�:b,M��}WG���M�Z�im���;�]K6	�ȭ4#|����m�d����Л�H�/1 ]��m�;;�c?T
VQ��D�s�:ڰ,�E�T��^,�'0����Ě����
>0,�q#��)J|ۣ�Mﺵ_>�3���}�I6�W*�s�|�5�S�m~Ew	��f�����Z����2�g#S)-�f�-2+9�*jz��O%��o��3��wڮ�#��V"l	� �JuU�8d��C��V�j��]�-�&�K(�SW,ը;ȥ����Cz&i�x��/A
���@Iᮝ��l��x�vˆ��r�d� �`�������o���8
��gFq��^��&%�o���9m��yޮ�t�#��G��8���p�9����*@Ŏ�{N�i��u^6�¢�[e�~x�-��
(�&/8�
��"�C�@��p��i��p�ȏ�~�^����]Q��ea�S7
c���ғ���H���K-
��<�]SDR�םV��KW�Qq뉖����R&��G5R��%��c'F(�g�i0t������`ag|8�����Q����Q��s�X�;��MS��~ΨQo{:�]� [�An�� �U�1~k� �?�x�t� C�p3�+�sU�"�;`�e���q�ߞb�te@�*���^�c�`�p%��3vz�!Gc�x(v���[	��s�@��j��R;7�ʈSs}%WU.��rʃt�{��Yt�:l�	k�^biw����b�:@�!�L�e#@Ag����٧���Ż�CP(� H(
O�YrP�Z2ؖ�Z�@��Q�*��,�:�`V	��G2u"�C��6j����$��� ��Ԇ�练���7@��!8�>�o��a~�����y��G@��m`y�[8�s��X��F���q$Щ��r\�5\����L��(��#���4*���zH�u��H�<����%��p��K��Zs�ke	�U{"�:�y�
�pN�F��V��58w�|8U�JD�sȼ�{��T�%��� }�*<��H�l(�P��w^*���qS�h��'�t�+��hRY�¼�]�!��6w�6*{&+�k��S��� wLn���a/����P�W�Hm1�Y���G��o�^;W;MRtO[(�nZrI@�[�\F8���>F��V��kܫ.�<����ӘE~~`2c��B6�)H���{�d��[��>��3�����_�,=TJ���QM���*�*]���B331��:ҕ���'�q*�����f��d�� �[=
Ӥ"QG���M(�7szs�/"��	���@7��R������x��'8x f��1�䖻�C��Կ�����A�{=�V��z\
�d����8!�8᧊m��3 H;��Ҍ��}I����>���ٍ�q���ѺR�k��IC�H�d7��ޥȈ��Ҹ0.���#f�0G�z��&�c����x>�4����Y5b�u�UqLù����.O�?`���O��DO����]"љ����L�����b��U�l���^� �:c�7EXa�\�+"� l%�cs����� ���¿�)2�6��BU��B�><᙭P�Z� 1s5���q��%���t�/�r@c�/�0L��}����g8�ݍ�	��1����M��_��uj��J��G䦬6��S��3��4��x���"1I����K��D��e�V�%8-�k�;?a5n���,9�7Q��M�+�Q���Ѷ��R^@7_CX������ߣx�q��K�8$2f�A�M��2����p���ř�7,�/f�"�`89E���v�6�m�r��,"r1��܏�Jʕ��W��o�3	P���K��c� EI���Ilx��ĕw��'һU�f��hM�;%��J�\n�W�D�@�D��E��*�y���;�U֞Ah��vc�u���7�̑9���Ɯ�>Ny5�2�ڮhCOc���f�\�i wF2D�~g�i(X�����Y�|xBJAq�>	rK��\,��5��_g����
�H����l��%�qPŲ��[iu�W�PԤg?M݌��k�q���`��yz�#�&Wssǩ���o��G#�.���F{iz�k��O��SMR�#��o"�A$��m�7�7Y�?��wɲ�x���x�~w������;h�>bNM&j�Lk-���#	��+��h�m9��-ף���廊yY�G���?������X�%��^S�`O���(�ʋ��ґƜ��C ��lM��o���4=�έ�|��}*��~ò�9~�Q%ζ�qp��q���}.8`\�q�\�㨩�����������;��VA�w��\�uTJ��ҷ������
�
)�)[���l@�4*��NH/���Dۂ�8�}P���5\>�3zTJ�GiT��zdAf \�M�gBN���ԟ��B�*G��<��S��z�q��A�{]ϕ��`��o���.�h�4�d;�/��"�Hډ�2��m}V>=����]�x6td�ka��tx�b������$���� �e���f���+PG8�)�?]%��r���М� _>�"�Pю	R݀� �e�j�}/ ��� �T�����1���e��fu�qS�V3�hQ<2K�b�N�����4ecz�+Tܷ�6��}=|�[��)� i3/Z�pı==%�N��e�ůMS��8GZ�} */����G5uء���]r
��m��;o'��]��ȹ�[��S;�G�!.�o��L��a�Rs큜���1>P�����t,c����@���$G��U�f�<�X<�ڋ薔���{�o��r�ԑQ��U'uxaˑ�kF]����1(�G�[��<RH�^AUb�CY���³��.��Gx�֞��7K:o�آ�|�9����xȥSPx^}�E��|ڞ��L��{7mm��k:y��+w��9��؃I�����l-�'_�Ʈ�T��۠4U�W,��)�t�KuAq�[�u��u�w'�Rw��Y&�Z>G�$&��ʖM������O��B�rϳ�Y��u����զ*<�@������0j,R0Mt^�>����H�_�9�҇��R��hqLӣ�����@���*���O#"��S��Pc�6b�J���>�>��f\HH>�)�ZG�F�'��S�✬�ΖW��,q��Bg��-��([8q�q�ob���[mv�ħЀ��K���WT��*{�̀lʉ���4pj4W�,��m�"2���k/S��f)��A7��xGK�!�j���xL$B�l�ʃ�m�F�fUhf$w8zz/|��q'mʞ���`'��.<�w��$|��g5g�p&��s;i;.s4�*W��W�[����V/$�{�k��5�FP]�N]�s K�bhn���!��/@9�Wh<�/�J#���J ��ED:$�K-˃^��B0����@��ד:UTO8PFe)��5¾�ݎ_F���>$�'a
Zٙd�̙1��x//ɭ��\�������^dQ��懢�ʏ�@d|�<���e���!/4U�P3���K�XL�.�q��Yv���Cs?VY/�K��ܣ̾p����xzK� �w>�}�aΊ�����k�-m)S@�\_��V*�gΗ;��<76w�u���~��{�+Ǌ6��^Tl����\���:�3�Y�?_�$�v�"���B�$d�ҫJYX��u-r�8��-"%��������!�)Rg�}���߃���*�����Ȱ :�2���%|���B�]���?��Hh�p6�q���G��P;�[�d�{�q�(+�և^Ĕ!p:ꭻmi� J���[�Q�Xs]\J=�2���F��+��A{��.��~���䰜�����9eU)��W�mJ��;��\�j@��P+^�5�R����<��o1�	�wT~�w���B���04�IS[��O�	#Ԇ�(dQ���'g� ��Ɓْ"���}(f��� ]��TM���������Us��_�v]��߉Tb�$Og�Ru"��Eۉ�(!Ƴˉ2{\#/�cS��ja��3�l�s�g`�Hc�#Ku��5�r�v� l/XД��٥�Hc+'�e#	Ŭ����H*���Z�-E4�\���f�����<<�Η�����k��\����"�rC2�Y�����~����p`[�P�����o�Sbw1-X"@Z������Ռ]��u֦�ߦ��͊}u��\�MQ��K`%ʽ�W>7�j�L��s$( H�8e)��UD�����8����Ş�FYΝ@����|�~IHe����Gx�ꛅg���%U%�T��JV��1�;�)7����-E������5np��	���$�@(��K�hp8�M�7�pH(��L��Fhn[��GD�\���D��^s��O?=�`L��>�rMwy�a�2�ic�.���$�3j�ғR��3��]퉫K�'d��4�y\p���R�0m��k�Q��1 +ںN�#u�`z0vf$YI�����Y�'�sd��$���ۢ�`)U�:R:x9����}���쭾����>.�,IP�9<AM���h�>̏ �����٪N�3^���U`y�Oo.�L݉�*R9D&�h�)PX�/�.�,�as$���q���a"l3\�&��5�ټ�S�:T�X[;I0459���*�WW�T�6�T���j�I]QU:B@�3������޾)A,�����g�9E��ͦ������g|R5�)
z�!%'b@�09(i&���0a����4 ɖI��K _����/U�&LJO��{O�.���+��9�o7��w���h{A̿�\U��!5�ʳ[F
:�LoQw�|�S^4+�EP�����ڎ��j���t����|�gY[N���ô7�Fs��2	;}z[FM�8욾D��CT�oPccЀ����4�e�����E��"��{�.���l#1[rlI��:b*x��;&��V9�x;�V��/=ԉPI�3	ܘR���/�u�Nb_�u�|
��ǐ�KQN#X�B�V�� Ս�FO���������{���xG�ٻ���+_���6�􃠍1�}Ѩ>�������_U��!"��b�fl�G���݁q�)8A�^����?6qZlR�P#��i�?6�V�L����j�C��
�P�&N �o;���!�X���fbX�:����D�GS�{�0� kV�t0"�J��db�ZՆD���˳������|�����ֲ+�r��c|Qt�D@f[�����3�]�r��8b��[���|�wa�U	~B�0�--O����\�&�T92�Ҡ�2�"��1U-�"2���i�?���l�jG�`=�#�C<᩿��9�V(g%*`h�*��pA8��N����.q ��K	�:�U�y�x��K�Aj�)U
�,���d-9ǅW�-]|�(w��[;a/'�sB�M��D?ZҮ����lF�D�r;��
�� ���_��1{�P�-��i���MI�ٷ��զ�8�UqV�v#2���n��F�o�D,)ᵪω&^�!{HYmT�@��`�Ly����.�1k��P,�I=OX���r!�z�j�2	���Stו���}���k����Q�I��-h\����
?�J����f�����6p��4��]�� �v(��[�s$/5�VZ	�����>�r�ռZdo<�� ���gl���
�ҎH���Ԓ�D�����-�b)Wά�0�;�#�U^ĪƯ��l�6����3~�m0,�'Z��QH5�չ�w��t��/�Tactyy@�"�Ӌ?s�4���GiFS: �J��S�c)��j�	4V]�B�:�Y��۲���nc�6�v �L���s��2k\���d�K�2�fץ����+���t�^�"��˘�d{z����6�$q��~@wPl�V�y�AeX����8	�P���/\���I���q��W_]�����&�fI6���M���[+t��I6��<�>o�r�ک���ĂBS��X�a�c.Z���CQ�5�m-�M��ɴ�ND�	�g�I�+P{�����p
$i!n�bU�� m���x�9.D+PO�p�n4#�ܑ�]G��(,{��m ��>F���8�`w��i�]�������7~ك��q�����IA�n�.����K����!3�F6ót6�л0֐�h�e��U��z�]�'\oJ>j�H��b/:
�|0�#���}�KC{*P�qȻY|/߰Y��������GՑFg"gH@6���ޛ�#�DD��%^%�ZF�GvnBRFD���2�T�'�5��= 9�"$H�
�H��Ƌ��>[���.O��WǸeŬ����<{+T1����N|���\����)�v��i0�h�0����M���/:,�'Ƣ߇A�]�����98q��2%�f�w�T}�/���Gq0<����/K��~VG�N�]E��
忯ھ��]��)�v��E����>� j���*�F���$x]�KM�l��
F͢�gf��S�������C�� ��wr��qţu���t�!t?(�W«c��%?�-�"��O���̦Ό�dK��!�֜�s:���P�B�8���:�2�T����|{]�����5�E^j�6$�s9���}I�ɲ�0�Z��<Q/ϛ�=ɢ��!�٧fEm��%�|Q�J��C�+�螋��UZ�=b�ُu ��G8����q%jq`�S��3*�/N��Rۀ%�ën���|k1f�Q� �A��9VPo*�Y�r���*���RJ�&%�50�%�މ�N�E�RB�0 ����oqW }&��z��rؐ	�UNh˖�QE4a���
�g�_E|���T�(����%%��/O6xHM]�o�.�A�᎞J-���EPh�=0�;�BiRf�*ʖ�vՏ⢌�	r\�����ت�x]��7�S����}b XS��)՗SC�̫� )��i���������#/Ϯ�[]v�R�"&�Q���l%��y\�+G���#K}�oY6��"kQ�����b�о�o�3e,�f�~`j4�����h����%t�eƘv� ��.��A��L�gPqg��$� �jQ�(]���9�Jm�&�3�#�֎P�C���ؾ5޺��Z��<�ԇn����b�94�_�b��6���f�������x���`���~R K�?^��Y�Xy�З
n�n����b���1,�A/ۺ� �`
��������T��z�Ê�޿��/���o�D��l)-~|�l�{�)�9�@߬�Q�b�i����f��o�����Ӯ��d���5]�E2�'�B� �4��GW1���A;���Ǽ�(����Mؾ��X:&���o�_����?޲� (}Ǉ�$��|b���r�(6nT;�=�����
�|XR_�ó�߸(Y��=�Fί�˛�h�{�m����D����~�֞�GL���+bRh�ݬ�M���'�Sh��%���6��"��[l�8d�C$��;h�"��1��[�w���7��+�ܯ"'hmLl�����⁨�a�s��#��-�/��xTi��ï8Y����g`��R� ��g*�Pռn���GÆ
�.��=�m��{�akJVߦ�{O=�ki��t�u���6͉��p��6N��?��dZ5{���H��!?�zh8�����&�&k�|�Ј��(0���ȫ~�A��	�{��U.�Su�=۲���

�+C	&`OߙzN%�t���ܿE�TO��8�� ܩT�H��VH�����J��~�g�����X�Ҝ�Lxd�7�pĥ��nd��pd|�F��Φ��w���0~�CZ�)��W��O�D\�'3�����J�%�8H�w)g�]�P�&���D���!a�EB�=>b�Sܴ��L1D;k{�p��N� +�_*��XcQf'y�S�I�]u+���E��Rƾ��_�˅ASX%��ٳu���Լ���8�I)Ͽ��YU�2X�a����U�Ha*Sv7��?<\=�%�˫����,�-Kz�b���2E��Y]�k���۾�=�G�E�XG�ͬ�v�����llFdg�� ��چ)'�*}Bd0�pE]#�׆���N��GB<����	�."�d����/�>9]��!�;���o����@�{��uK�w�r��P��e,C5bY�A|�C��tH4ǳa�p��jv�n�	c� Kɶs������E���T����%��e�~�aò&z ���k�W/#\%YU���W�Maq�"r��E�cNgt~�{���������	�u�9ZE4�q���`�ذ��	�f�'�l쭙9|�o(���y'��s S��/�i9���)O���u�F�}�axa63���S�H���_5|}����Lh\0WdJB����ߏ6`����|OLX{�Om|�����4?m�'I�3A�.��^*?��KS��PXW�4�HT�i���j�?�n�]=9�b#��>����b���b��b�0�Pv�>'��c}�W�?Y�L�;�£v��\S��-0���dp��!�ͺ8v��_b���!ۿ�@ ���׳R>�!y-��g��yD٤G��ؾYn�0�Lf]'�,F�@��������9�`��}{���r�9[Z1�q�C�����6��@f��s�	Ѳ�LT7>�4�GS\$X\���2����M�
D�Ņ��r����(�NU1����Ρ!��~�M�]b�+����ЯmujJ���e|�cy�K3��t�F@�1�V��m��C�Ɓ���-|��g���8z�E��P���I���%Z�sm�c&| y!h04V͌��1Z��㉓U��:b;�.����*��>f��xsɣ�mv�1Iԯ���t�
�h�1��"#b� ��KA����������������H�3.�h^ângI�\+����l܇�1�/	"�+���V�_�_�)���B�q�l����(ү��+�m6�����V�[oG� w�B�z�!aP0s� �>2*d𳫋چ�h}�
�=t��sG`#�k7KU�����=�bLos���\4�@��Wb����jw������jl}�Ѕ蠖6�)@�x��T)���?�6�}]�)�ް�Ys*z�	n���P��y��z���%	XUh憾Іmԛ�%b:1&R���`iӦL,��|%���42|e����Gk-�%����ѮoH��[x�6����[S���B�j��9��1[c��_��$���N\�ܵK~�u���֦��T�.����%��oû�º��5w�Q1ݏ�����8:��`���zĕnQ��Ii@rt��wk\��2��/���m���=�e��R@���x2����	V��+_�Fs�v;?!;��O�x��B�<�/r��R�~:x�L�g�j�І�b_����{�� ~��a8��5$�L�N>��?�z�k�z��~8-7��%iS��$l�ܟ���3�A��F�*m�Wt�g0i	|��RuH�*��;̄�o�Ň]?�T�s�R<�XAW�ncK��	F��0"�#䪎�ؕ}P�M��e��IH{���a��N#�ļpuR�y�;�!����*���2���0Y/r�)A��L��<�r��tI�֙��F�Ҏ;<��&r*:��5�r�͑� ܠm�n��Z���"e�-l��j�,��6[e���[����{�G琙w r�aG"���k+�:Eg�?�ؑd���<I�'��мg\�l�&���.���ߊ�U���n�|�j��K87��J�gMH_^hƎR��SC�\�bb��*���cO�F��4b�Axm���l,8����;cWM��q�*1A-���Ǜ�P���ҁ�����zi��|IM'������5����:��"�)�4�ۄ[u����dVge�`, ������Ԏ����l��i��Fd��<]��|!m!>��ϧ&��p>��M�j����C���}���QǷR����=!����@�)���h�i�"TL������4�w��։rU	>�Y��h$�2�ɶO�j�zen��qEz{�L�s����̱��u�X�J��Z�B�z�'Xԛ���@"U�[��Zo7�z	�O�V<L|�*bl@5����.�=v�h��z�b���5��������>l�(����S�~+^ٛ_��xJ+��r�;"���0�O
\(<؊��>m|�MZ��Fy�w��HsI�*��=�y� c��� Y��C)���^�_H�E$Eg�Y�SN�<L�pk�e�9���t���T?m�I���s��l�V\��P1�!1�E�(������#�1�K��hz�.��� ��Ʀ����vB_��J����L���6p9/� �j���/��e��i8MQ����˛�ŭ�����c,ۓ}�(�ɧ���.��}�l&��Q@X=���e��M���o��]9��Fa�S�#�ǽ���g��H��10;X�K|�>��)O�s�g6.�B�"�>�����Ә��a���ȡL�dfEB��"ڌ�KON� r/�;Ք3�����&��$P;�" �/��=�a�6�x� x=$U~�&��!P�x�fd4"��`<��"�\��Q�%���_O�
q*�e�m�Y��P��T]?wr�ڙM��2	0?N��x*n�.�y}��-y�������H-f�������7���KD^3�@]Em�l��\e�gn?=��	���z�� ����Z>��ç[X�F%�n���'!��>T�u4��,:G�Pد�k&���CPt�Oؾ�߅}��%k���$��:��v���E!�b�cn�C����]�̻WQ4sDK��4k��,J��Z����/��zd��Ӣ������=��j)(�R6��M#�յ��E���W�g�ֱB<2�z��Ď����4s�`v,t̑~WsA�cuF�.h3��]�wY� �.�y����#Z}Ef�<*k��Z���N��TΔq;#D�|9ܣ�R�� D�{��'�E�I�~��m����{sv�dƗ��`��ގ���_�cTh�r,�4=���w���!�u\�͏gPd��7RU#9̺eK�Gg�|�R��lu�	�eǗ��@Dl���o��^�+�)��+�v�~��wLX��d���>�zL≰��G��TD袭��4�8���lj ����7�j����~�(�n��/��0�V�C\��+��_�%�pTs[��
b��*�g��3�3�t����4����z��w�A�ww��2�n�M{õ�n�#;���߬�֘ �I��5-�V�ɋ&1s����k=r�%��f]\D���̩�?Yr�
 ���f�Dx��+=�?���B2+��s78�O��?����sֳ�e� ���7��SV�ɿV$����@�>� a룅�Aq����8KF��Q��s9nhMW�}�s��ݛ�����Ǧ�P(�*e��d ߮�����I��օ#u���>�<�p�)�澹�n�=~fh��
�`��?O�.���"r�����"X��F��>w9y�D������W���%�u4x�8^5������#PW�l6��LM�y�|Zq�ݝȬ2��P���|�L�ŵ/�OW���	C�H���K�yt���'����hÀ)~� V��`d�
*Ǳ�f����Pz���1A�ih�I���t�Pr�]���?�']���w�F���2mvg�?G]��2eAu�y�D�Y՗��hkt�z��!�:����$��;�� ���:�S���iF����rh�,�hs�N�k&������`�\���o�ee����1�O�HQ6�_����_5e�m�aU�q�GՐ^�9	�R���嗧�5ٱ�~�#�"�o���M���l�ۤ��;XdE-����v~E!���0�bc՝v��`ͨ�g���3IO����S�P����,�:�w.�u������5�e;_	RW��,����\�T�@M���!��j2����h�U�}U����B �W�'�k}�@;� �O�����6GL���Z�1^��/$���I2�R�菛�"�%��MQ>K��oSb���|Ek���M鑭�W�$�&
Z�?v�R�����᜞2	n�DY���ɛ�i��g\Q�*r>3W��o��!����(q��$�ǭ��3_���/\%#Rw��W��Jg$Tp6uq���I�LӋ�q2V� ���c�{�:b0�Czg���4����&�H��p��Nb
Y�T�f�����w� �=�����9�e7��  ��.��<$8[���r��3��� ��r���2@�m����Q�v������3P�`hZ//2a�L���������P)65i��M�܉�! �Z�`������ ����,�hG���5]��i�j"s_�����ы�.��c2���B��涝�K��9�>�����Ҭ�Jx�f�Ɛ<C�k���p���l�Aϑ#�V����;�m&�mQ����YK������m#��1%3�~5�%�6�X�	��d���ܽ-�"XD��C������M_�V*i�7-~�z�������]�]@_��x��۽��I�(�}Ƭ��):����
4�M]�جA�E�K�((�-��qL]E�QcZ��a���D?�S� +i�#��Q���t����J�w>�����ޚ�h�� �|oH��B��P�blԕe?�yW�ŗt�ݸ��O u��\�� %# �71ӛ�2;K����i>���^�99�����	(�E +0�WJ�a'R��������L9�.v-ک6��<��i:�]��N�H��ի�?ų4\x���r�_@�d����֣�|Us�c���<��4z!Nhe����N�cq����B��Q���L7�d��dY�7�V\k+<�X��'�J�V��ytS�	���1Y�j��Yt����4?���S���~��/3�^
@�;g��[`��B
i�!'_PrI����=ٻ8羱/��MY�)ͥ^<h��yL�M?�*�~+a�=���#ߣ(��T��!S�:��@p���!{g�sT5�Pn7;(�gU�1ׯ{�G��״������is))e+>+SW��/�q��U�a��-��=��� �k�S%q�����<�t���	��,�jDe�GPg�g��#"�K�����"�U$S.��%���ڑ���g��Yc~x���&��R��UbG�u��ґ.}��r������-vK8�-�)a�+)�\j_�,�r�&_D��#���5�xρTKxq��(�d�4����E��݌*�=�L4�X���m�M�f܆�_iQ����S\�\h>�(4:� ��؆���Np7�f�NևA�`O*Bu�R�l�p1V�,��?�3Hܤ��_ g8��?�m	p���_��ty3��_f\���zG�hI��XG(�-���!�|Qh�9(�f �p�DC��}�|�CW�� b��G�)Y?
J
B���G����?~�;���d&�VCK�3��̐�I����5���P-t.���[�ᝧ���l�����KB_��:8d'�A�oϑ~>8��1��n���c�5��+K�$\yu�)b���cxǫ�`�-c"�Gos]@1D�7"��\g�(4�U&A�L0i
7|mBym�^���lQ�<��� yӏ��@�^��s���_\�w
#�Xzas~g �����\,)`���z�l�D�w�N�i'U!�9��='�Gh�*��gLnӾ8��>��M8T��^�_ՆP�w���u�ϲA^��%,�-̵V7'��^����HZ�0�ۭ�a�sYLyM�o�Xחz��.��^H�s��>_YJ�#��S����H�c��A
��4����� �V���Ϩ,X�m��l��1�=�=���FY�{o����͂廤Z�+����s��6@��۷ni�DO�1ТF��	h���gH{�U�
2
	[Qæy�� g&�/�q�оd�����鯀��OS�!��{�%��zC��"*Rb��"<�C��!�D�y C��x_��r�:��°��oez�B#�� }�ٙρ�E2�7�[goq����i	����&�!*���B�ƻWϽ��4v�>ê����*�5��Eh �+�Y]~�°A0c	�/JFU&��S0�L9�g�l��l����㡧��#�/G?�{I���Dg�L��gu���Q
�w��DB�����6��cy:^�4�����{Mq]>�T���.8�p�C��<�'B#%v���[J,��6�|����K��`&_&}Q$�����l2�*2{Q�Յ��U�FBHB�ԩ��i�Mq^,��"�䰱^�'�J��r�>9���wϞ}� �w��Ql�t����.RJI����uv�#yy�>�f���ŵ7Ы��R����nW�3��"�e	���Qý��_{b9�ŕ7�0�37�k���x{q��<4Ҩ��S�N1G�>Ny��d��2��Ë��LT��Қ���O�k���Ue�����JY���qp�f��(��sS�QB"H��!?�����*!|@t�tT�߈���Q@����t�pc�����wBGe\}����@ �\+��ē��X����8��Y4 ��l;,#�O5;�Ph-��En���>�z{�y��EOh!�吲���j�Ġr���p�y�'���z8�9��++ڝ+B7�z~�5�qW��"��.��D��A^)/�D��ד�+-���HLtYT'�ŋH$-_I��λ�=�mYr.g��#�t�@+�f����01M. rF j�pA^���Xi$6� �X�RT�W�6�t���q���p�-*��h_tY��X]�[J�y`�ɥ��P��Y���GX�TI����.�ԼZDa�H>����M���P��<$[xZGV?���:ؙr�K���fD�YX�~41N�Ƶ&}��0�	�Ą �� ����x�w=?i�mf@EF���3�I�cq��#(�o9[�8��>U�0~�Z:0��x�W>١��������,9�S�D��.���z��7�Q�u�fs���� ��oe"YCaajj��N�9QL�Ԯ��B	0~�%�KGCȯ;� G���.CK��I1���u�x�V#��>]�Z�!L���?�ƠF�M~,ؑ�ed���\��l�s�i���+�)E����U-���x�UV�9_��b���.e��>U��ag���f��!S}��
ۮrC���6��Y�n�E� o$��r�� ).V���&8'fn��>dK�J��L�q%(m(����;gn8؇��l��͟)��[�]�~	����Pr�=G�jU����(��<�C#Y�O=��+>��+��mC�p��}%�E塭A��[���/ޥ���,/��m�#��nL��:��)��hױ�l��nþ����2Ğ���2�9���0w���J-}�p~�F�9Vw֠O*Ev�����5�'�F78�2i�F4�.s�⛙��8�;���*��t�O%D?v�7{��0yOt��	j�D]tn>���u��䜕e[�R��@�e�[�H"yҊ�|G3�P��Nc2���:(\�/���42�߭rzQw�^�aM�� �%�����}��e��P�,��Z%��Gݯ.�?�O�BҁFt����UZ�d�]�FED�{w��,�P��s�J�H�S�Mf��I� �t|�=@�в�Jh?d�
(�4���"�gcJ}��Yn�kĽ0�C
9\z��l�-�<�'�q�5�֨k����#���6Mc�l��� m�׭��8��G+L�0�8ԙ]���u�vk�+�s~(�~�2O����)�~=��A�M����w��C.�@a�kqn��g��Y�F_ y��F.����7LhJ�J��!���C#A�J�e�L8��f����ɀȖ~*Bf�����."��8�~��Z0R�| j�y�^�}y�v~�{�bq7��8�����F �d=&��]�2���3:J���=�̯�W�m]ǵd�wJ	�Wet�Z0"i��J:���5�鎌&� ��o�I�RF޵c#!�X�fJ8���H�(�B���%�W
EvVc�T�z����>h���_��D7R�A�%�W$����qj�+wh��bi�U �����\�Ù�C�=ؚ�t��?1�9���q��i(�O�#�(f`�3��[&ˣP~����.��0Ƥ��\�i���t���W�<Ny�V������V(���!�+,��m��,�PD�~�����%�]��0�3kq�o��-��ާ)\Jxm[��>xJ�0N��s��}+�JKZ�������!�v*��}����ڿ�����i��I�Ps��5��=�ˡ��p劆���pj�EJ�Ṭ:�����B����5z.<
���eK�PM���/�Mӄ����D�it�=���E(��S�h����Z�:�#��'�D!.i��S��T�F�Nk��CZ� 2$�g�ؤl��+lLr��-�����4�%.<����Cǎ�>Ds{|q��Њ�R����Fla5[��v:h�\d�?������#㏟es_Sdu��~��O2h�7-q�<����!o�mz�Tr&c�ȳ��,���M�
�_cW-h�D��F>@�+����5'	[6�3�2�7����+���֊�)�^ԏ8�X�	(׵��ԜF�4�������ԫ�9o]d2�4���-�}�����O�P=���r���TR0�����o��r�s8{Y��;h���ܒe���j�����^t�:T�d~�'kjֹ��Dl�:$$�e;��._R����ՙ��O!|j�]��z}M8B�0Y��h��?:[�v��*��&���]��b�I#+p(����(xj4}ÀJ�i;��m��'G��?����/���5�u��G�f���y�[B�zz�P͏���}��b�
l^īl�{9���PC��;5�Y����5�P��C�t_�/�ٶ��S\��'`�U�.��YѢ��nl��+���_e'��Wx �_?&"J��#�e��
3(==�fǥ��k؞��1O����L��k^�������!�I��+)��ߓ��CV�8�Utw�Gq��b�'{�:mwy����T뇪�M�M4Zg�S�뛴S��Ԧ�n]�	��ju�P�w��+���i4��=�sֻ��6�!�Z@ ���sjf����
1%%�G�¤�>�� ݊�MRA��L�|5�e��L���)Z�(I"�X�ɩ�6U`��J�v���#�!�@�,H���Ym���_�k�$�  ��D#�H1���2 mNiv��|	��6�gy[o�Ic���J�C�_��*ퟯM6��u2��L9{q�L���~��Hi��$Eg�B
����K*%�a�`e�y���	��R�<�ft]�~򾴻�����mA�@��{GhԶ�f���f�i��Ϛ;��ܴ�>,���6k]��F�(�õ&�~�H2m�%l5��5�=�粴y���ާ01N�^��ގX�oV���SC�q�H$�5��w�����k ���2��$���
���;:}��s����BD�j�0�
_`�t;,u�*�H�u��T������m��w�9fk��<M��Xi���1�[�1����1���:W�K���/v��*@u�*>��Dh� ���$��=W���uz���P�v��?���l�_C��Q&&yӏ�k\�D)���]�����;y�Z�d$H;�0�_b���$Ŧ����Q��WC���s�p!Z:������k҂��%w��B�.���i�AZw��L� Z�B����;)��U�i�*hz���f���W3�,�[j/�#�+�[4�L�Q��D���	�ć�f/@/�9����
��g��dE�]]��n'h��
�r�8��K���PL�w�>��/ �5�����C���n��I�<�o�)[?�كP:�{`d�q�����T�����L\)!���`�\�܁�]t������_�sE�|�.8ؼ>�h�xQ~����S�����#�@������u�n��4�v2�L�/�So�)���yo�%�3��p-H�3����I�褡�Yz�$ߴL��ԫ�Y��O���7�"��o!`*�4��_����*��n�b��"[���g�U�;��Ƃaȝ#��+���t?jy`�pJ�8�T]�������9^ΓA��rJ���3�_�8A��)��osx��]��qkm� ����)7S��,/�H%=С6�7��Z�8�R����H?���z�R���KI�|�� Lח� �)ƀu�k�j�V����M'{Tۥ��� �tI��@�a�Y{�2��~3}ծI֙2���:C�S�굓�#��AY�4ZĞ=pTQ�$��B3������ٚ@�6+K��d!�&���u��\p�d�S�x얛~�gD����e���X�3�
-�.���{�l	�mk��0XSO�*@��aY6gޥ2)�o����</]o���}�]s^�xQ��V)`��_u;�yfT-���}��nPԅ����~r���1��ֽ^��?�g�$6U���d��A�Z�Uϵ�!5ɟ��Rڱ��3(�>A!h�Y�L�>k���E.��26FI��0ZE�H|4npet��͆�i�+��H^�Z1WY`��O�p��.�'3�`��w��%I2]�4��Z����~x�!:z7�����8�Y����*r����	og��RDv�n&p���!
�Q/�Y:BPS�J x������������1����_�y���_U	tä���X��M�_YC<nNZ� $�.$��ZR�q�ܲT�!�M4���B��]�Y��=�nwIl�fCZ=�k͋\�w\b.���D����cy�V�v*�$�W+C�
w,bbjG}�M��9�t0�&�� ����$�'���ek�{���N�O�l�.N�%qQ�Ȟ�U�	c��b^4�CA�����\9 ?�0(wox�؎��Ib(��I��gb�4���ͨ��s�ڮS���I^eq�k��m��H��]�4t�2ں���c� lQk��,��?�1d�	{�~�u����x��X�TF�a�馘g�۪o�S=2���*�^��j8�yBU��P)�rJ��ь!ܨ�������Uڑ��.��A�ƄIw�]��Ŧg[k��p3x�It���W7V�ĸ�n�DV�����n�$�-�s�Q<.ջ۸>����P7mW���9rD#�����h���77,iC���7��צ�1Eä#�b��|S"Ȕ�_ox0��j��C�,��Eg� 0��md��<���޽���H	�[>E5�v/�I�}��"�T�=~M�^SѼ�U��:�nn�9�̀-b����p���Ӂ}\���H�~���M�wy��'P�x]3�I:ԧ��l��$�{tD4e�}�O�������ɿ3{H��l}�d�*c1���w'	��pS�YH������E'MB2h�S~Jk�kU6ySz�Nr�m]LQ��a�,$랻������C���1
��g/�C����n
�� ��Ȓc�R�2�_S���\`�o�W��"E�4�)�x.�k0�߷��{� ����~�H*{���cu����Uo� �-
��9�2��ܲ7�9�0��߃{'a�g�$����R�e^��rz���Yp�Џ�T�iKeځ>i�
U'-��e~���4��su~C���ڰ8[!t5�յ$.8R�X�<Nvz�g��4��r��MOx�D�ֽd���a��n���:f��D  He��lK��"7p�[q<~ ɧ�0����B��v1Q���(�.3:A'�澁�2�4vȦ�C֎�w��v��_Y�#e0��u�����x�{_s��Ai�����I��U���� <p���9u���s�l�����c���\i�`(�]^��جâ��($
J�
ĀWB9�j�*����8����yt���_{���,��(eyحc�������!n`=�茉��5�h4/�X��x��%f�f��EB��tm�.�f�ãF$��?����b�����k�����	��K�N�� h�ǥ���4�2�;�1��C���E���l��/ɍ���hC�_�YZ&�.��أ���D�!����C�	>-�ЗIZk�o�V�.o��K�[|j���D�[/�Pt&ߠ�x���6�N�Ci�fT$�<<�F[*2K��kl�oo�&���j�m�����ε+����g	!��-��(�&�%���8z�[��p�~��I���3����|}�5d>P��?���� �h��6ʟ�-\v����0Q�Ҏ*�n+t�
�@�Y������ʑX�)��'�Ձ� geoj�uk��m�O�3��Y��լ6��,C2ȸi<�� T���Cԯ���, ݼXZ�!z�Gt��0���:!K0��5����dZ��t��4ɸU`�������I���>n��l��zoS8 @�~�K��|>v�kZ=��Lv?:�I?�)�4<9����ܺ�,l /{v����	-������f��T��i*Q ��}4R��c�O�1��L�5(y����޵1��ڢ����扺�+���
WxW $0F^���7A����|M��[��������"�f���Tz�9S1 +�h��)��]Òq�0����Dֈr����9���Yw��\P���`\s�/��G/�#�;�!�t�s(��D�+�?��q�)��NLҖ���2�W7�]c���w>WiXޝQ��P��)�!��?�|䯟%�����Gz�����l4Un������Ie���K������ג�G��T�i�?8^.̽�3h?0i�m�؇�=�@�e}]$|�(�gg�����
��D'�u�,������{��U����J��jJ^�[�����Q�1%O�+�)s����dMA��#�X1R�"q ���n�˖�% ־��1�޵�냥K�b��^v_���N����:�/e���� SA����b̏W�v��B�SZ��%��g�������#�)�Wo�Eo��v��04�+�/�}B#k��3U0��ڢ�,@�P�܋�Z|Ԑ�׼���JҬ�VO~f!�G�:����1!Ͷp�ӎ��J��[q"a
f�B弅6�]h�y?�G�������ҭ؊Q~`l'˩UҀs��8G��g$��Lv%/��2���E�`��S&���*��<8T��gv0�E��az2�ǆ�>>c�t"�^�����<�;'�<�}���Z���;C*������>R�J�=˜ ���V�݊+=XN��.;�^$��>+����P�q��b�`z���Fxw7�4��k��:¤�P�{�ʗ������E�G뛠F��y>~��J-úk'X%(Y�J���S	DCP�*��8�i��ʚj�֞����p�n��8�P<���R�Y�w�x5��\��i͚%���6/�Q�ђ���ـ����E`s�M��4���;ϑU}L6��/���D�	����G����\�9�a�e؇���7���w}���n�`�x�L/��N���Tv[�B��W=V���?y�N���j6�M[�m�����b����l�N���4�3�N�0�#�fPO�HJ�T���ͫh8?E���rtA��OW
0ڤ�VۙY֤�,v�"��F����@��rF\�'q��l9���C��YA;�iU�J�drgtE0���j��3G�G^���M�/��|UJ���@��|vG��M._ȭ�~yx+��yh�~��yd�3v���QI�ʈ7VJ*����o��;�1^�Ϧ�eF�O�v�iN�(�)�}{����׋�kWh�V:��r�ٳ�u��$�'�U�_
�t�$��T�l�]Z�7��V�'�"�j�H�k����Y�.���8q�T����1��F� ق��c�!��Zo��SC��}�� �P��"�4F�)%�Z�� ��h0>�\~��N�UsJ�4q�5�֏�ə����s��}����c�
i��El|9��?:�� �"���F�M���+��Q���׆_�����\{S���.p���,�l���]U-T1J�	��C�)�qJ����bP~9�	�<Ǚ���X���������$����-ޖ�s�~������ь��<��L��Ct=�7�|�h���x-����nPA�#~���~Y�%�Z���ÝԱ�<r��s��R���Г��W���K�%�?EW+TcY����>i$��ǈ�MSI�v\NE��ƜT�˖�ܲs�M��qᚺ�@�
!"��$�ѾB���t�`�Uc�K� ^b'�A�1�����F�������NZ��6P.L3뵃2����ޏT�lXZ?�=��b[˸��Pp�T?�htG6�3N��)��Ζzݵ�?�η/5���l�@��X��y<���l��C1�u�*��r�K�jbx�ilUO���/�3��gh��{����J��\�L���ô��Chүe;���jWɁ#��w^��K\崾��_�_�\���渵�ӎ�[7�#Y4vNm�]￠-�ZNm,�hf$1^_	F�ˇ�q_�\; l����X�D#U�miӞ���
T?'��0�o
�EJD�5df�������pP�E��:`DMy�� �� i�mi�LX���@%������I�s/H^Ru�������f#�5>��l~c��1��1����SV�>f�MFj�,�O>������ۊ��6D�r���o��U�L��wQ�V�WK����[l	�����؃%T�d�B�Ѷ?��vXvҌB��U{�0���h��SJ�N�����Ch�z�\:���f�D�o"�y$�:�*��x�#�W�4��P�ɢ�94��;�wu�	�`�Sv��4�Pg�#5)�|t@�yf�	u�dnZ5}��)�{�O+D�W�Y~�_��[��F|�>q&�	z{�n �G��oMk+��>�[�ì8���f�����}
-=y]�=*�?�{4��l�oB��x'�ܯər/c���
>�(���Re�ZJ����耷�Y�D��U�Od\�^z���'m�:�6oVqP��g�8w{e_+���V��-���@K��Ƚ}w�w�uO�)��H`5�L�D�0c	%/��K�dN�Q����h�:7�9O��a��o��½X[^��$N0aEӫɢ�3�U���]6MC���T�z\�=�x�Y��K���-&�E[JN9��ן�9�%q���p�}��~t��v��t�*�z�7r�B2��u?'��3�� �`�0�1��h|�7r*�x��e�	����z����$��SGA�S:`_δ>	ā��3��]��U��S�h˔0�_ k��8'k�_��`�|��չ}���^6�Y�~�S)�t��)���4y��nָ�#Hf {�f`�^c1�^4��^�ޭ>HW"��8#��@`��i���~󟀼�%�+�����wTҪP-E�`,���6&�d�Uj���`��	���������3`�>�F�#��Z�޵��������6c&M�󤢳z���4	(�o���]���Ҋ��c�Jg��C��o����ʋ��L�`�뢑�?`�/N�IEl{�� ���w�{�b�d��5'4 ���	�����������)���2C:�%��ɝF��Sl܍" Wf�ߴ�:7�6Xk�#�,�/� �y�$V��?=H:Ԍ�U�mk
���c�m)�`v�L�ӣp��`i��nq�Q�������uUT�TB�|Ѧ�+O���yG��7��é�b��3p9�PyCFG��5�A��D��������D9oS9��)\�V�~�ꙝ�,�|P��|.��.%O��F���������$�q8ñ4E�Uf3O�v�8̝���hR��e�����+��?J�ո��g�t�J	�R���S��#W����`b:��Ŕ]�����GO� 	�9�~����"� ����NU�74����:�J��WI�\�k����h���٠ b�іa��˟����+��ed��l�prf�6<�VX܈���������6~�Z�t��"~ީ��vY1���^��!#
�@G�wo�I��;���i�c�w�R<5X����a�I:�{�1�}�֟��ϻ�!���8g'�q�NɳN<��M7�����Q��ֈ֌����C>P�(�y�f1�T��T�:�B[�JZ��WSa����p^��/�~dw-.���DU�g�G]�w�a�-6y�R�	��Q�e�y�m���0FM6�b��\�WOd���}	SM�0�I�R}��5�y�yA��b�c��_�����X:t�<v،}�1�T�G^C����������J�@�B�!�w�� C�(�YZ�a�����+��I�<��ِ2.� ��zJ�����a��Y����d7�Q`	4�����wx����'X�B��:ƃu�c�ᖓ��b ���l�����4i7�ǉ��c�SQ����W���;/�(����({z�ӫ]W!�����11g��ǋ�_�F�q_��A����C�s(��We���9��sQ������:2N�
���oH5.~(��@%2$:	�{���aW*#���#�QL�\x������y�.��cv�F26��K�ȴ���l��Z,A%fi���&��!ǚ���h��<Ί��u���H/���w���>�>i��J>�Ǝ�2��� �5~Uu&v!�j�d�7\"�\���;EL��Ѐƿ��L�Z��D�n�j��%�Ի�M��n.kcY�x~��#
��@�W�� a���l��#-`B�:5-�C���Z�sT��:��,�ie<��|�Wva��x�c���m�	q9���R�4�dG.���롺Q��H,z/���X�����Jȱ��6Ku��a�'Շw_A_�xݴ��V7W��8��� ɟFbKt/�F��bǀ$�e��q���q�<A��q�4��1gC�}������M��!� o��
�m�O�3*1H�dE��lP�\Q&T��% ����Bz��"p�q!m�q=����A��Z7�1�t��Wb�hPn,}��
����ӆ��-�55~X��U��A��X���26�������s�S��q#�ˢ�H�j�A;Z��G��΋s��x�C�w��e��<U�ʎZ�Y�5��#5*�<�ô���سw_!�K�{$Lv�B�wz��%�t��zlh�b3o�IC?%W�/��kUN�2�Ĝ�h�O�W��ώ�<���í�ƣul{�Ld�sK���\����w�j�
�ll�w�AZ���7���t(���MߍfDM��p|he�z���SY��.��T�/#}��v~��%�Y��]c=c!R�D�EHܒ�to�'���N_;u��nE�-�5A+�X��?WSw���~f=R<��,�8~U]H갚�x����=b#w�Iesa{�9�ԣ�)���7Q"�`���s:�f_γ��Yؽ�Ҥ����[��e �sd�Bs�)^�
N����t�}t�b5P།ڰ�r�
��`oϒԛ'z���LPGU y�@���7���$��ڛ{��L��n��ܒ/`��P�qN����ZU����h&y+(^�@������*攦8��S* ����o;���=�R���� ���+}]��ݼ�V�� � �b0z�!������߼���!�hۧP�8�HQ�N�ر{��T���B��"b۪��ܶԢPL�|!��vg������$i+vȭ��7�	銮(�eÀ�"I:�}qD��9�,��*���I薤MY�	��.���)\>'����!:��Nz�=�Jv^Ё:^[+M�ە=ipl*?4R����H��;�V�y�`��(	55Ғ��;�+����}N-(@Y�L��)۰sq��}6z�_mY�Rٴ����:�J�-b�n�rf�F&����ҭ��@Z�\@u����,��sz�� �����Pb��m�q7���V�i�lE���T%<������V2�FRBF�9N���+�s��T��^�e��I3�������t��	�c0vН3k�_�[	���b�R}PxS餋16�{FpOD@B���S�QUȊ�+��i>�3[�w��l`m���:8�.���h2x����)c>��(62�J��lH�9�\�ٓ�������/Ʋ헰 E������a��=���ؘ0�p2����=�^:t,���?���W���l�Dӱ/���ԕ�D�{JfEU�	~s��3��eZ�|����#}�E�ǫ�pBg} �I���B:K�����bd�i(t���K+)ݛ��="rENTI��A�j�n.��FQ8�ZfG�m�3���o���/����Ui#�D 1!�ΤO��]�K�"z�D<�Cҷk��0:H�p�q�X����G-�D��b �3��J��$s��l�U)�(�$�8|�զh>��S�E3��w�T�m���&�U�]��FԚ�eb�xUNK|�N�4�2�6ݽ¬���F՗�
�-'!{,g�ZC(ƭȤ]��OK�2֛q�Qj�����A�U��g\����gU�4ס��
O/D��N�p��q�\��ZY-��(߈c�tl��/P��;��k�s�a�vH�ӂ�}���Њ��o��!�}�)�V���'�HAb�M�z����jstc�XÉ�^x<<D[x+�kN/k���q�`����y��-������Nb��J!MO�Xǆ�^%��0�ُD�-��<v��R��H��	c_,���IJ0bS9]j̾�@��H5��Ug4t�wW~cU�fo]����CT5Y��R�2NF٘�U`gi���o+��T,���ŇE���K} _��n?���m�H@��,�p_8��u����[��\��Z{�S�|ҡ�B �L/e|��k4�p�g<�M�E�U�ʒ��Gi_l,���c��,�G���W|:�gT"���Ӫ�?Kߨv��b�P��j2�ݦn{�,���	HIh��������g��lfH�
�d���lz�6ŕW�j!0�fy�H��r>#ش]��A�o������4H�W7S(�ɡc<D�ć��4�\����C˦��q�?b�"��Z�� ���{�37.�j�RU��S�^Ԑ� р[���c�l<Cչ[�z��.yW�J�z��5S�=�P��C.��s遮6�O p�|e�J8UI��-�!�0P}���_��kew��Sw�T��/*���$�Hk/r��8L�[A��$�~��ĭ���%�xIhL���Â�)s����v��;Ks�2�H'j�¨�H&Ir���1����o�Ō��03h/�W�۔|L��U8tm��fƫM�0�E"�4�����I�=\ɉ���`�N��.�?/r܉��׀�����'���'�-خ�� :Oq"ci��B��8����3�4d�����=A9��{�j�w�D�N3�� ��_�*kPz�
���M >����$ǻ���$RXడ�+9)]�����)4'�t��(#�a���;Y��ZŞw� �]�Ԃ�`�!��{��l��9�I���:H��(�/�b���=�UO+2U�i�wWk�$�����t-�����:�aXD��U>��$`���3�i��Uɔ���c���Zy�k���n���Q2�~�Pˉ�7���j������=�ک~�K��
�
�>���Ĵ? k3=�����M����\������lb5�����.����Ѱ�-��3��~5ܴ�K�u�/O�az��� ���a>�ǕK:������ �9��|((�+�H��M��|H�#�e����*ns%�Jz���&F<?�
4��߬Bz�i�"�ָ������i4���3ɂTf$]N\%��$�%��{p���67(߄(�m[�;x�
@�Vh�H��_����ܩҕ��y� t���c�+*U��6$�q�j�-q[����� ,�6�'?6d�0�s��U_�4Ws�J�q�����e�:j����s�k�Ż
'����dN_	f%��A�U��aMI!��<�.$}_���8�)W/�[e�e�Z���SÓ�)���;i�"���i|��&��<iZ��6�x�9�P�!7��b�|�O}}P��FǱPwJ&K�����j���s�>A��Rn�v��l
-a��M�����o�FA!|wTy���{=MI���S�!援bAͥC�q�,0��J�a� �<�q�&����vY����Viusx�ȇ�q��K�����m�-�a�H��1Nʗ�(lu�|7X(���IN9봵�~�(�e��ވB�<����ĸE{��8�'U�:�e�ĭ(�πT�+1����+TS~g_釷���L��0��F�\��K��S���.V�/{$�8}�rݺZ�K��1Æ�zUL��<я�Y
��k$@uZ�"U2���s�Ż�nϮ�!/֭T����p�����z#�e��p�=u#��#�j��� �&K����&9�8�DIG���W������} ����+(�������r@�ex�~y_6v����2�����f}S#��K[� 6hI#T��i�vʭ�A���nD{�X���j�+7<���*�z�:9�����D���Y�ˡ!���<������nQ#f�)��+�&6$��U���/�]X�~(� ��;�rLv�3i�ڔ�ߗVs½h� ������7ݱ���$��'��{���O��wy�Y���
_�sv�Hs�Z~z����"e ���Ȗ�K+�y�L�A�D[P�l$x���a?���gM�,X�8�iN�l]�c�@��:ӭ�%��ϼ{Q(!ܞeDM9�~Rh$m�:f��qCI
�(���8��]q�)����ٝcђ�~|,oì^�Ԇ%��(��l��7x�R��|�V�ȶ��`VlƃF��^�� ��_�I�����c&[�`����a���Q�w	�!ux.�?Y��S����*�LF%v&�4'7��"�J6�N˰�8
"������Ϡ*;]�_�Y�� r�D(�1zz;M�y=ڃ�_�6/�̩��n|@�������E��`��/Q��%=��D��Hdn]c��q=���~P�pqL�wQIG���H_�w*�cZvsj��?`Uҳ���t�����[9Q���k;��h�0���z�;�b��Z�����?�w�$@
gL�}�f*��,���������ۧhJؕ+IJ5�B|�4#"�ͼ�����	P�P��y�?�%���j�� ���E�:��L�_��J���/J�c�k�ɖ}K~]����q�.�EebO����T�ȯ�a�r�o7VhF��S���e���a�B�\N��5��(����O���m�f�ËR҅��<��P&��ƌ�iH�S����h�<�:�P����L���7t�E�p�9�W��:b���f]�A��5@E�BѠԴ���Zފ�r?��և�4��-{�$kdv�@Y�%�y�B�v�F�d0ќ�Q(�F-�w6��k�­���'��맗�H�r�c���xmO ��' ��pM���M΃Y`ۘߋ�q��V6�wD��(lT�Td&f$�8�>�S4:���q��Q���1KM`BY�X��.���m$tWc�����/$��.ߤ�)��2���V��c���N!��@~�6z�b�崁r�m�>υ�\���f�7*^s@�s���*��'���jؕ\c259��wdÜ~m#��&Ϡ�j���S�W���:����3�*�-0���[Y��cD����7�r��_�x����S_�;P��rwڞ\T����]�d+��8���#h��I�ދ<�4��� |�Z隯�x�OVƪ�:o��ĳ�ԧ�$���-Q��{Ɋ�F���6���e'7�L���,��Z�Po� u��Y�)[[,�f�@D+����}�D��i�Q�aW���d�Bpܜ����N,f(�	����u-��Ӫ�}fʳ{�:{Fd?��OP����w�֮ӕxJJ bN�U��{ �%<w�o ��_���((v�J�=ED7����oK�6�anfuϱ�B�jIqt���H�ЮԦ��z稼?ð樍��@���2����.\�٥�S��2��]=Y+��R��yVE!a�c�y<نjك�+�#��!<cY}Uw�y23Vm*�r�u��"���y�p����r�G�{yxT)�;n���W"@��������!�cT����m��B�V\,��N�ܡ9��pW�`�����r0��1Zc�ڻ�� ����j�L(*����� ?��x�X�E��^�'�>(���!BO�����}���L��=	i�*�fPQ�]_�Q�
]FCV� a�qX��3D�^_��x�J�����+���@_^�y������0�N�]��Z&wBH��:��A���.���&Њ!�KJ�{�3H�\��[;�����zs�oD�3�HGV�	�u�a�d�)�? F>���iM����IR��Lxf��#��[pá9�A����Q�O�4���/<W3��]��M�[��_iA|�bG�-\Y����*��>��߰������ޚ����,��V^��#�E�k_I��1�>�X\�c]"��"�MH�ǒ	�Cb��⪥�=�5�2h5�p�6�EbcC��M��8|�#uv{ �[�\,�a�i�|��i�X?��'���գ���I_��F~���
����jB�y�����'�{��	���E�,fp=����z�G�S9
h}p�_�&.'�8�oU���ɝ��绢��cxFE$�X�Y��W������0�J@��~��#ո&HB���I��[S��I�*�@�GR)3�Dn�M칛��
+�-�m�
�Q���HK�r��&ԟ�	d�UD�ᴖ�M��!G�m3�6�O�2:���Zx�-�R�0W�+�L`[?;Y6YԬPز�n�|�6$��[��"��C}84�Zc���Q<��?
D������nU~�Z�� ����{�3���Kq�1��Su�T��FtH�͔z�LcC��� �m�����2b�#�F��.��_�h4���4�퇵�+��1��
��*�/
���ְ�����i�P_�"n-�e�]@m	m�f�j�F+��X�?�����l�K��
t��d���ie���Fo���o~��`%��B��~5:z�i�T��̘�����ovH/�9����y���SI��<W�I����+7#!vkP�L1G��Ĺ΂v�b8隭���ɧ�����Z`���������)�L\_��ơ(��lbAB��.����>m��7���0P��A���L�y.��勐&�����=�j��֞'M;Q��@�(���88&뽵rZ5f���`t��{{$5蘋!k�o�  �C�{�R�}3�y��.�C�5xN�U�6�|#ѠdW`�aϩ�m(#�*�{�@��X\�6�]��U:	�|�k���{�(-%V"�O\���O��:j3-�p���n��_��08�C�����S'�)d�u� �^�_�C�R1���o�,�7���.ZB~M�)���i�@�a��V�w�5ooǴMs"^0�𰾉ի����xg�:�k
!��g̞��H2`�2��ZB�6j�"�b�J\Fa0�����('7��FIJ�CMX�6��A>�J�0��~�g���Ϙ���Vi\��2U�+0�����@���晊�PѢ���n�nC����:��R�Hy�D&&��`�sS��O���a��D����w�ح1!�8����*8���ԝw�r����C��}h��S���yyl i3U�|q�)�E�h3W����;\�u��]�m��$����īv<�Q����yeI�:�9f1�}�� e)��B�qL�&,�Jt�����o@��+Y��~λM�����U;�<G��D�;�A���P����Ĥ?�ž�u�~vƯa��f�oy���?�`t��h%��F����B4o�㚆V���(.��FO%6�j͖�7W(�E��w�*�vj�R}e�O�[a�-O5:m�p��\A`Y����0�`݆Vy.����tvɚ5,�-�oH���S�<"&��0f�'�v���x�O�$�uR�lN���sQ�Ҡ�q �+~��Y��U�G�1ĳ�@�^qK�Ԏ�`Ϸ�C�'�@p�8@���'T���n.��_<��p*��'C��J�Z�[,<E��	ҏ@�󉞏��۫�D��H���_�m��N�P[=2����Iע�R.\�X%�R�`�9%"lO�Z$kM���d
�(>/ޜd�i8���z��nֶ�Y�n+1�����C!��0����G�[�J�㣨����}݆��*�n	�T�=�;(��\�;O,}[�AH>j �1O�\B)�t�Qa�)���D�ԿV;v
q��:x�u��8���9��(��Bf����q!o�)n�1��"�t.���sO��l�!(�p����̫��j�P����k0e �m���3b�<ɚ��V�O�F
�"��/��Fx/��(���p9���Ƣ#�6%��Dr`n=!��#��?P�����%�-q��v���Zؾ�/W��8��)m��DJf���&k�
Ċ�Ƅ���ƶ���bu�N��G�j����� ^B�ڲP@NC	��.�1���W"i+[%k���[);�
�4����h�t.���iY��̀#��Θ�W�D�(+U^$�I��yt�O���]��\�[k�?L2�/�Z�G�'���e�w,�I�H3����.�;��(p����&66!�;���4�2��RƵ��� �y6`p/(������+NoC,ԉrI�.s<%(���JpZ������Ӕ����eb����'MGd|���"*��1Un%�=�Э��_?�ILc�/��g��d�+h��e;���3���X����z���G���!Oq<R>`L�5��XI� ���lg�qQ)>�^u��u$�ɾE�����:����#���������	�����,����)�R��5�q&���ӓ�b�
}��_RsD��g7�3?>\�?P��y��s����������j�N"(��}8�
���6NͻI�7b��'�R��`��2��t�_���ϭ'
��c��F��S/��3P_t+v���2�"��o���v���p�_�!%�j�K8������'2�պY>��A��֨��dR��Wj &�l��,&���[ܶuq�0����N��C�*�C�뼕�C�n'��U<u~��XL/���L�^!9kӂ�Su�wŏ����U��ZۍC���;���=�Y7�VXk�]��7x�)d̀����U��YP�ӑ!�(�+�Bި�C}��E>'�h��N��'����ۚoD���O����b?�Mx ��.!��يrO�������V����9"1iwqN��@oz��b��m=Ą�,:<�l0U�#���P9|q$+>	9�~%%�|���+�:�N�x�1|d.��S�0�
ē�Xd�VHGpyg���u[{%>y�ըQ�_���S�b_�؊��_��T�Ck�#�;�[�F��4�;G�/W��G�m������a��k�{��4�v%���kH�[��e�l���;<Y
;��V���?����W[��'�,��K�siY��@a�|���q6� ��R�p���v8FkЙ� �o���xg��H����C$8q3�ZW�	

r���ǰ�r�q���(I�ۉ�HSAfcr�i)� Y߄���ɡOo�c�S�2%V���<y_:h@AX�ďs@�(��V�~6?ny��!��dB5�Ƒ���q'��A\��1�N�<�✧����n7���H�	��Y_Ѧ�6��t���5��ym��Ke���c���l��Q2b8W��I���fV��8��.�\����6j�w���Q�V|�\ħ�D(+�!���I�ha�N�s�霚n����&��>b�~���� �����K���Qd�����q6^��X	�H1���NA��5�JsYx����`���k2��h����g�w�hg@�C�+L�E��>�a�/mC��S��%���o� ]�4[��ud�!����8 	/��+4��D/n�|CpLŷ�o��o��C�'8���l�s�-p��yu/'	�&��"h�_��ZB5��<����-�O�����˸xtl�w�}�}i��ڼ�a��i���o�2�`��pA_��>���Y!L65�IP�Qg8�Z`��rS��C�J���`S�Ң���Y�C���BP�{G���RJd�WZB5j&���f�������� �A�GA�≅LB�G��ꨲ�g�j��hc�wZM��G�m��8��0��"���1��`e�������"I1^��7>��έ���P]�Aoo()�.��g�L[��\�!s{�3ŭ,�@g5�G��	w&�!���&_�<���ʬ�P<��?_1Tc/gM�y��r�d�%	9@j�g�Z�yӍ���f���ǙHʻ���m{���2ޒ;�ò5�Rz,n��5L�I&��kln�Sk>��f(���.���;ױ�*��ȵ�3��`لHd]�+N��cЌ��O\�@"�),���r�Գ�3.{O-&8'l]^��{@N��������&L�,{��)nB��'8��Z?��Gǧ�p�sL�8�Pek��Zc�m9$�N�J�$#���PO}h_��):C^$��ِjuݤ(Uw`� ��	o�
rc�S�C������m����⁗�����w��#BI�[a{�^ �?\Hb<@ΰ��'?���c���\fǾ�&Pc����[���
K��S�R�"B:@�&�����b�&�U�h����y"E5��;8!��q4�*K�08�ϲ�*g1��f���p�\sx&jr��3�8��/�/� ҧ��\O�p��|3l$�hsqzQ�Y]�Pz n��`�1ς��K��fK��P���Y4��w7�ߋ���q*�d�S�1&�Z�Ѐ-�r��*Z����"�C͜�=#%�C�VH�� ���%`H,����'"�h?r��>�O"��A8|УH�pL@�����?�i��xׂILv�� �%K��T�WRF��O�7�K�3��'��qGʨ9�ݝ�qF�LH��U��m�$-~<���;/e�0H���b�?	J9,��c��I.Wo�f�LG��9|e��-�?�6���"Kn�C!{V�t���Gp�a�@.6�L^P�?}I%�Q@W-��X��`�~òON�������GA���G.�f���24�*AVgw5"����s���>�	�Z��l��z*y�6��w�_�mV�	��b�F��Kl|AMnbg����uG��dŀ�?9;�EyL��8�ؘ�z��������{Xި�ƊYNw�q��ބ��#z�m�����3�k��#f��B�7S��O����#��8�����9vU�]D���^�p[4��2��r�N5�R��S�gŐ"Ƚ�9�~Q_���*߂�<�OGDv�/d-�!Ikb��y��&ךHY�����yg��s�ߊB÷D<e~ɑ�I�SZ���-E��Y�Zq��,����i�9�nZ�����]��WT���Γ�����+\�0��D?@�,���m��܊�	<�7� ��+d�I�=���-��A[�PX����r�2$LWq����9���2����-�,�+Z�a���k���^�	0�r�J�S�`���cq��@jl�~-�V
ߜ��U�Q6nZwc��!�}%E;[�������2��r� `�~+|ҕ10��������B�ȴ�B|K_��r��W=^�F@&F��Jk
|-��[�s�>�!5!Uh�>�´��|?<A����� 0�vs�՘��qS�a"&>�d�e�o�viVI���> ���؀8����Qf{]�-p��F  FȒ�!�&����́p�+_I��f:�3:۱͆ձu1�Zcf��8!A��:�����X�F �����v�[u?Wf!��+�$�Qk�N+��M�v����{)}���y�����ׇ�wn��j����IC9`�ǌ��-�$�ܘx{-7u�"�nu ����<�~?��.,l����E�ƛ��U�A;&�'���}=�8�ˁ�N�1�$ z`�N���3��=gx~����[K~�d�T. `��CS�o�&�l٤�����
�O�>==�llDW���cT�1��	;��*�;u-h��NS�����E�oU��?���=T���g��an�	�;d�xT�D��H�A½�qE�nM29@��,�������?!�rT����A;^߹�O��N��O%�o���4���� �s��
I�{V�!����W(�v����ET`���I���~R^� P�#Qd��8"4p��}.˪�R���Ef(�/����8�K,��Y��H4UBc�O����N�A�(�Y�ñ�г
���5���8�ԕ��E����<��t�,������ܙ_f��y*s��@�J��%E�?WªTC���]7{>m�[ʆ��)p�S��*y<t��o�����]��VGC��~s�X�3j���ϵ������t`��ME]P#�c�U�XV�0[��8�����l	�M1z��š��(�<�I%&PB����j `_���AIS�~'>���)nXK��M�Y0:���J�^��7�N��k�y-���B�FZɷc	�|LD��:�p�rS�yn������ۈz���n���8W�P�2�^&�>�!�����3\#�n��{�WU�}CrO��l��q��&/�8�d�r��3'���o|�NE�΅:�K�OI]�ϑᴨ$�eo(���W(�2��N=<6�>�Uy�G��D��3n�l~f�h-�j�-�(���y�J��k������т�r4�J��J��?�� 0�{���}� �UQO~�x0�][�Xa�=�~���c�	��g�V,c��L%�qk�#������V�@�Ư��V�O5X3N���ո�2�������E�7�J�6gnŃϭ8h��8�7�i��'o�nZ�"ʽ�~L�L��1��s������;kIĮj�~�rfZ�EjY��Y��Q��h"��9Y	�~����5޽@���ωA����ʛ� ��o���L7oy��9�c��/
�b��l�!*�o��?� ��a�=�d�d٧��hhݟ�Â2�Z����1��̞B��Q�.��e���6��bp��W(*�O1�<�f�JY
��P�Ԝ�6��'3E����s�~@���,��Q0%6���b)vy}u�JP���4G�v1���AȲxS����~9���6mS2:/���r~�V��r.9q]�6�S^>@�Ə��7S��Ỗ�*��6z��2�עX�N��紩�J�t��U�I�*a�g"[ �-��c�[���H��ҙo� ��7j k��ئ ��ܳ��T�hgd"���G�vL�|�
�k:���9��f� tٰ�WF�A�|�{;�Y���B��{���{���U
�Wkk.�jG�H��D1�^�� �����f�A�>+[߹��������u�$�F�3�#���t�m�#�a��fY��3��=��F�^����I}%���%KM���r�o����2�H*@W�`D5M-��t�V�_" Ӟ��vl�yQ?�pNV��N%{��x���yfRT�ᔕK���r�^��u���s��s)?����C!3��3�H���.�i����hǴ��'�y�_N~��{d�#�b�t~`�!��ÿK��
�e(|���������c�ؿ���F�Z���}���:!�z2D�ip�ӵ��H,�q�aǩ%��J����Vjw�6;� �z���*�d��X
q�[m���%�^��H��[C[�}��\���jf���\S�(ED;�*�<d��Q���>�=�	���b��|w�03��ra������j��]'o��u6E�'ܾI�����"m��B>q�MG/6D��o5��v<��Q�BZ�@�7�G/��IQ:,|�e.ɡ�<3π��g�,0�
Al�G'jָ���XPݣ@H۾�z�.=��J`5��2�	7���\I��Qꜜh�$�<�Dk~����>)�5[N�~zT��)�����$�Ɏ�v��+��>����/��V��DO�T(�%���8�^��.�pA�4,͇��鴤[�K�����z���feъg	�~FǓ���q��LAb������n7;,��me�d���+Q�h�Q:���%�e�ey��{�=%t;p�R>��S�u���Ƶ�X���:��hT��㇉��L���~�3T+���䁧��b���!��5�|�MNu���A��5I� `n��b��n��m
aE��#�S���$�x27����6� ~x���òle{<nMv�}Æ��`U�sΫ�t��S-�m��@F��)������czK`���o�uQ�+!�17�Ћo׈g)b!m��6��Ĕ��]���B�@/����M$/F ��`�����<���?��K�=ĝ�Dč y]l|�9��9���dC�����'�L���>�f�!8�`�{��o�_)u�c�U�U�oם{��jV�Ɨc�p��Da��ۅr��^�����&���FM[�g?΢+���w�i%V@?���bZh��a�̼�n�+��L�F4��z�s���f� ��+m��ɫ=Q���A/C
���[�|LG��.Z`bv((B�\��i��2}�C��~48=I�X���p�C�D��m��y>�/j₋<�Q��`���m�
�3^!���HTk�}�}��8��\3|m��H6� $ָ_bz��e�~Z� ~�=�/��̏�e�Y�,��3!�/����⨘��KF��MV�{��_%ϲ���A����(F;�>��X�ָ#���C�Y���]~ ��2��s.ϡjw	_FΛ�g�-�8�F/<h<:��� ��Z�97���^<X�X��J��F�N
pD�4��Vr{�Q��>�O��c�!T��ֳ��\��yc�)�o�]��9�5S/2�Jp���._> ��9Y����K>�v8_O���9h��3b��8X�2s��H�1��ۦ�'�J�A+��<D�	&̟���R��(5�c0l4#��r�ۤ���:�ϼ��F]H�ְ�PZN
�R2M-!�j�W���0��w�
u�ģ$�ɀ��\���Ps۴HӚG���B�;� G�y�����$���^�X����A	Dv�h)=��@�D�n�k�cuEo�q|͍�3S�SB�5�%�pD���h�D�0S�J�|\�LP�2�����+���C�����ݡv"�&/e=����xE� -x]�7/m����V��������@+�n;��9�  �J�,г��!$y�R@�f����\�'(ݸҟ�l�3RK9!N���)��K*Y��RgQ�PzϚOh��$�b]G�`�p������3����'�G�$�X���!��Bc0VX�h[eG��q́<m�0\�{�I�r�ͺ���`�|��n;sL��000iHr�
�����a�B�0f�z֫V%8?ux��M~�5PvSU+8d�q�6���_�q��۩_]�"9`�=�;�%5LNNҞY=1(�qh�~p7b��M�Y�f�h��ݛ����EρC�K�I��o���#��g��2��%8vʊ1z^�渿.�U[�,��AV�G���z2�	�����=�O i[�ءL���J���B�J-4D|�U��K�d���@QH�H�5	P���k���>�7b(|�4^s����5q $KYL�� �u���$�.���W6��QeP����Ҟ�"���^�@S��'��0H�FaϞR�i�3���h����@���������ǎ�� S����(I� �[^�`:Pq������G M7m�F<+�b;zMPq���D  E-�u��U�e�KK� 	e��R
X�� ���[�r<_5�'D"C\����Eݮ�y�5�B�xӘ[��!B��;6�C�7Ab�~eU;/�G��K1}����<�i�� ��)vweV`T��mH��TR�V��	i�&A�Ru�g��:~Ǫ��&�wY9�7�ݻ�^��A4�����G���+E��bz3u�z�sP�x�"�D�  �4�(��~�;��#u��w��8�v���9]���	(h0$ς���P��*����>���y=���z�md��a>B��ǚP���.�w3M��_�:sL^��R�V�_F�|��I#��=XB� �����s��?6/E�ƓZaq��.ٖ�e��v�����6/�>��P�_ �m�ԦY�jN�#���\�1���U~��[�;1�۱�g�/E����f�����Y	�H��B�;�<���^�����y�I������ �c���^Kf}����B�_��ʠ��V�Xrk��↕�j]p�3k@P����@K![/�+�~�
�n��}������(_�}=1�O?!(K�q��(Z@���ʁ�*�iL�C��ǢV��E�����sz�/���BS؊6m���� ;f��JB�%D�*y}^��au�$pF�/]A�wLKd���eA�?7�Y?�/�14b��K0�Uȼ�3��?\�I<��7������
��a�ro�B��x���;����T���ʟ�X���'����(�/#O9�����A�����vj�g���������D�M`�ͽ�'C�^c�oz�.Q�񓼯Ju6�Wn/�0���W|�lY�)_4Խ�����	w�#�8�z9���<J�_cZ_tU�1���p�~x�qC��|�/����Z([N�%J}Q xyzk;��/q)���7~HYBhbG��7	t�9��<)�wG*Cr~e~�GZK3���<Su��I�X��G�=��F�Ƅ5] ���J���9'�����y�\����t�C{X"�+�a5����Ga�����	7�ؙ�S~��`�]��q���b�XS�1e�Ijk��0[��]Ͱ�(�z�+iFE����|�{��c�,���Ll�"�=Z����c:�����[��_u�������1$�Ӯ�� �e�T����əNr��paq4@�Ү�����=L&h�S����*m���ClT���`�\o& 5]�}c#�7R������Iv���(�^�'��?��EoU����"�Z�͊�Qk���9_�I�c�%��T!���;/Ho���k�p����4����$���ۻ�+����8��?��Ti��]��io��:��������jT�/���OG3޼uI����#��W�!)3�9�Q=5:�T��\�����(K8M����\Y��kLz=���g�<�N٬eS�o��;'{t�޴��K�~nW���q �x ���8>F)�H��g�ג/�Z��	.�f��߽�d?��GG���Y����� !�UA�L�a�z�����	 ����wo�֙:{PsmGN�M��my�AVZ��i �N�T�ɰ�6��zK�U9[N�\��>3H;��D���̽{�	q�oH�m�[ʞ� {��V2�vD�>b��Y��g�{0X��bT��Tj��@c��hJb��OӭiXA�#�W;wD2������2�Mv�0 ���\d޽o���ka �w�>t9�#��^0���M����@��H��D��.c��@>�#�"���B�L��e�X1၀w���ݳ�-���:|-U���By��{��ٟl
Q��tY��1�0�b�������t@tX�>�P(���+-�U�����
rױɒjs���n�={�ZB�2�Z��V���`���֪�9IS���f���N�0!rp��W�I�/P��!�9�8Ad��T���R�� y��҂�p�G��h)���ZWË�W�%<���u+K���5�u�yѮ���E��gn
�~��%/	�s�h���
����?F���Ul?�=z�?	����Į x4D�k��3�������|����5Z�GYGb,Q������L���zA�X�i�|��]�	�J�,��8����I]�;����G���Jf�U�^������$�DHoh��hF��X<��%�����o^r���x/�?�,�"ֿ�~�;��[���w�)(.l�:�x�u�~���N��8�%X%�WC��������62�J�R��d����!9ղ�&��[G��܂�J:�i�|�a�*�2�Z�L� a=�	����+y��|��|�����(��/3]��qg/�^���yr�83��1;1��X,�����C�7O��e(�[�^3á�A�>s>G����yulA~��z�W
�b�0턀�{�䤳��,�ca���rg�A���U��}�����C�l�Sk�1M���8���lQd����Z��~���ʟ�?Ki�~��Y�a�H���@#>���7���$,����٩ِ� ?�^��֪S���@ NN��VN_ 'B�w�K�'���<b�7�Lsf�B�T�)�G�Eu���dfw`y&�K!��=Nl~`y��h=�Z�kE����R���H�N�ǌ�rIHj[ߗ�^��]�Iv�-���?v\���������@�G���.�@��'Ķ��9	̽�4a��	Ł������Z�� `�3B����d
��U�"��*	Uz�M��	� ʹ���I;\aFt)4E�� ��$0�i���A�i�*T�͎��&<��%i' Cm�g���`ǧ�@N����>�9T@�+s�|N>k5?Eq����1�e�e�=���u{pm 0H*�H1מ�u�kK�B����ޙ�u]�'Q*?Z�Z9��¢�� ů�EɊ�9$���;�׈�&���?�|sS����d>�u�%�I�%���C�4�rX�$Ó6�h*�S�����ٰ�~�ǡj��񿾜���3}������Ȃ�Y�WR�������/��ɴ��9Y?��Gp�-��~M�ŋ!�~�>/�D�  �b� �@90}��5&dQC���${S����^bwzEjW�i��A�����A%�ߛ�`�T�6�!�1�s�j<ҝ숄ۿ�y" P�Ԡދe�J�8� _�{�sZ��ػ��8�l>)���HZ����J�W��6Q�*iqS�)S(�28�p��=i������U���5��\7�w7 ��1��;_ۤ�3�����>�V�?�O�\�tV�/�����6���Ҷ������&���T���Y�7v-n��H-6�
B��d��f���.�,�^-8z��k[��9^_v�$�-�?�lNj�������.-���K�4������c��,�������J�aB��ҟQ���
�)[����cw��<.�]ۜS�@��]$��)��tI�r.�+׾�R<IYN&��l��ݡi����j���&���Q�GI�mD������ʤGTz��b��zi�?��b_�E����Ӏ��:�M�y&�B4Vso�W���O��%���4��ۭ�|����4$��ce9&z�J�y�(mؕM�,�������#�����Hk�G�&�X�ێ/���@Ƃ��1�EؐnH�A?Mz��X1�!���[PP��[�(��k#�m`
�`+�|����,%@D�V���yl�#4S��=+�l�nZ0jU���l�#����`���8.�>��~�EM�6� %g?h ��/���+Mz��� jޙc��*����qC�4$:_�1�Q�B���Ql9M5D�Į�>�����_�4�S'��|3���7؄悾l�jx�T�H�H�T
����y�2�we��\3T1���v��2����T(+��v��*:�S�d�[���D|�ٷ >x^Rԣ�M��H�D�n��SJJU�hq���TP"o�
�찺�C�}�(OQ[Ӏ��k�O�B_A`~'=�P�υ��| H��V@�&�xpX�/"@F�`�kM�&��6�����羮��/�Z�;��P����6�@�ܫ-T:փF��t.�4��p4S6I����t�	!_��T'klvw�N����;�k#���{������H��"'��)5(�@���/pwM��<����tik��<2ڦ�Vj4����ƾ t�oUXl�H���Q�0��V�x.1�Uld슷|T�����JP۱��%7E2�0��p��v^�J�ȣ[4ڴ�O�o��tR�z$�5x C�Dz[�?�4�`\��L;�{��Z�Uҕ�Ʒ��804;�����4|9rMZ�u7��DzN�)�֒P���D�7��d�kQS�^ࢉ}�S�u #3�k� ���FGs���R�ꌤc�=E���(VrA'�Xd˱��~���U )����x��"Y=���!�HϞ�ν?oU�
Rg�4����瞦��mO�����&�Z�� �'C)Q�%,���.fQ�Q{�:�dY�.���Y��"���px���;��s�����"��-O��q�A�{o~�P0�=.�v2T\R:g��Z�[􋇭�����\��h�uI��Jh|��T0�3K��
��[EK43���|��u��r!B�+�~��#7�8Fl�>�A�ߣ��O���*�Nꥏ�hh�֫4f�e	j;}B�#�?�m\�kE�&�F?P�S ��-�1��J��N�����η��33|{�^K������uI=��2�u�'�4�у?%�,�&!��oڙ#��	+��-�!�n!Ywc|�}���&���J�Hk�`=B/�4�!�OCz"�����"�mZo��k�� ����><}����/�	�Kn�1ނ@�g��6�=�&�N��Ǜ��Ar��k�:S���R�S$�Lgw�U�����^Ao�u�p���n��d��t'���?��YQ�E�>�T�L��n-��e�rG���9��>��-�PB�}r
�wmԞT�P�����ŵ�Q��t�z�t<��P�:P����Lt�F����f��G`g��V��/�6�,�t:b�Ki6��"n���L-�䈷��F?�b<L^�F�g��_������g4���c��.�<Ͻ/b��A��J4Z�}�<*0�b�����T�8$ �_`�C-�K�>�EŗS�i ��-��n^�5�$8,gasm|Y�1�,Hf��8�5{��Ź�"�ֽ��X�/h�Z�p����Wu�d�b�@vR���'���P��'"q ��)�C�`��6����@�@��!��m�Il4�?>���������A��` �}�>a)�Z���"��1�hyB���X|��y�A�y�Q��`ha��W!^�b�%��%+������Tm-O�)�~�#~����Z�N�^׶��7؂E�b_�����UW6��7��On��}N}�_u{zɚ��
gg[�til2|�Q�������s�2�e�G~d�A(?��s�NMS�{t�CS빗� Z���� ���J�Q��_@������%mz�h��l�\�;���6ߘQ��n���Yw�Eږ�iM��z�h��R�� Њp����r�!��~@0�:�8X���is'��@��:s0$�.���*x\*�y���P�Q�s�K2�W�O�f�uf��<�i�2��J�uW����[Ü.Gl2���g�vw	&m����	�� v���z2C�j�qIL�M�HU�^�`x�/:��}W?�ׇlWQ�_튢�Vs"�&����0�Juf�5UYˍ�?�H��9�Q�n�ſ��{:M�¨�-,�Sm�VL���u��������6��7:1�P�m� ŀ��z�3��)4��
^
�� 	B�q[X�@����Y��i�VӅSZ*E�X��Yiyy�P�f>��p�5�:��B��� �=D��M�'{bA�<�I2��P|��Ϯ��@D�t��ܛ���7��~`t������)���<�6�� �N(�%o%�ƣS�=H���R���A^�"������4+WN(h�����;�YvCT��R ���&�n"H 1��0U��mO�_�p&���p��X�IDI�(�H��e�!���|0�!y�ׄG\�ΏHa��T{�Pޢr�v&�{̣�L�>kjJN�:N�l���bݶM�������r�/�F
5΍ŋ�3�t�Xl�܇g�H��� <F��.{�M�uՎ���ʂ �����#Jt��)�w����D|��w��)�V]�.+Z�x�ΤS�����&�uu!���������t�tuZ�N�/X%��������L!��v�(��
��YKq��%̧woT��vw�L"�Z?x�(���s~ۥ�����p:�ı��W jշX/+_��"�!1]�f& �kʣ��W�Q0fu�m��%��3�3/-��Sc�64\��|Ж���G��Ki�%�lr!�crj*ڵ�Ok�y��T�f>{B���6aQbQ&��su3I3���X�C�`���A ܲ\������N: +��s�챏�?
��QĄ��`h��v����M���bꭗ�MǐNz���`ٌ6����~� ,���-ݹސ�J�����?B��]A����p���S#Y<�46�]�W�n���_�8�S�|]�Z�C�����}�:-?g)=}2�u���TF&ޚ��
>�V�~̐�b����M��3q@}J؃9�R�܇�z�xT�-�+!�#30=��V�����+�,m��8ZOB���k�N��S�_~��M7!0�w_�c|v�L��rgq���Uؖ�"S�����.{7Mx?��nz�To6��^r	�y ��N�^� �aV�j�w����R������/_mh'���������0U�����{~oŌ$�ɰT�a�ߌ�?���7�+Z�e�]3$��'\3������V�2��ޑ##�|#�U��q,̦=��X1��]X��x�"�
e�b�͒���
���1ei��uD]�y�n}�Q[����s�L����c� dJ�Ɯ��u۫����sH)U����'�Ѫ�e�0P�rUJ�v����(8vs��|�Y���/SUa������omWs���@g�(lF���E1:<��C
!��$�u� u���>L�O3��\� ��J�F�V������k*��k�)s�hz���h�_`���}�eE� b��n���w�LB�΋^x��[{�`M����O�E1F3K������3V�zK�3�h�	��F6����W?��k��{�Ơ
�j-��m�]`��d�Z�H�ýc*#���:^�Q&9S$�҉�6�p�h+���J���Vo�oK�8Ҡ�;��h�Z3#��
����tw�������a�2��2
�դ���V�M��� Μ`��$���7�*��1����`�=����̏,zј�sSߓ5�f�E/t��h����pW��<q +􇁂0k����=�+T���?���˙�S�+_���#/�m��~�'��nUm�mqć�9�I�� ��+s+X{���0ot��}:t��4������@������#L<ٔEUk;�>Ѣ`��w�oT�Bǝ�w��lrd.ޏxk�#�CI���Гԩ���vB�*AM����<��4�����=�
$Z��<�ϋ�ӊBPj�:t�����Ǔuhg�4F�7(|(�7���& ���d�[\ɵ-��5:9�C�H�.4�.��T���M�3P$7[Y��t'B��v�
ß[Z�k���o�����F�9��~
`IAF5�u�!~\�;=��}�ZP�	V"?�*0J��|�E�����~�
����I��q8Y�A��<ﳏ\��y�m�$A�!���͠O�!�\I���J8@�86a�!�]D�a�Jڥ ��\d�eM��2X�3�,���l��F���%	�:��[g�1HD�{���EZ#}����8��<�$jF��*r�+�.�o2����*���d�w��e.�<u�^�
��
Sk�@U�z\V�@W�`����oš,�ED}0�7�g�����]M�U�(!�{���RʘK]ڥ!��w�����̃?������|��2N��5|�[p�9<^&ݻ�&xU�=�놜Yw� T���TCˉ5\z�����b~� ɏY(�����O�2�e:����n�O?fxEA��!:L-7���JjC�$�/�%W�gu7Ǽ��mm�[�{���y����FpH��^4���s�����������Ԛu�rz�A�S��ag�j�Y�-�F����(:��p�'�qL�)�b���qk�k5���T�|�=ʱ1�������:�1���h�q��� %��}%D�u��M�X֜01d�)��
Z�#]�-���<2,��Ka1����4�"����W_C;`�cDS����������ٗ��b��&�:�^�I���2S(]�A���&�������]��ԕ���R_">M����6���G��쪏�q�&o*�x1�q��B.��R[C5�8I�{z�b͹7�7�h,rT���_� �����S�ڊ�9�ؖ(="�<(!��Rp�(����V*����gjD�R����c\�k:ͱx�K�o�w�bx��tZ&��n�����pZ�lw^I;��*�dZ���@���S��)jOPd+"h$7�z��,v��β�j��j3��~�pd^ �D�W����jl5�T��6�\
��/���"jgJuO��i��p��9ʪt�)zj�^�㵇;_o���\4��[�ڶ���C��a*���&.\$e�Lm4w������v��|�a1twFE-A�-�p6�mW?�S�<�d�an:=N�UR�(��y�nw�L�d��%��6�� H��%�� R#���-b���N��Ӈ��ۼ�Y#�َ��|�b4�c޳M��/����&���6�M~�V�%�75
��w3�'۱�wL`�t2��7ܮ�x�٫����0�/)��|������5Ȼ�3�C���{��̑�<*�}��u���U�����³�ߗKU�*Dm|$���Ia'#�òW�e���D�Ks<�_E	�#�6�H�F]P�_ճeÉM��	D4�	�-�@e�[���8x�`<I�֒h��˧|I�5�����TO��h�	T��͉�'W%��߄/��F	`-����k�x�k���]���`�}M��o5K�!�i�6{J7`���>�G���W�Bs�����O��g��Z,����$�( ��j� �p	8�Zu(1��&�$¼����!ȣ�`�Kq��؛=W��e0���Û�E#�u�*����J⭓�T�;��O��j�����H����A�A0!&Ӟa������`��lz;�ٿ��E;?WB��%�ݗ�W�Kk��S�p��~�m�M5¶M��*�{h�����l�0!�h.�-�CQ�Z���U�yZ��ql�YQ?6d�C�q�ߨ�I��z�Ӆ~Y�T5��5���Ș���}���jfZ���~����e�el̓*q�A}�7vWP��b�Q��h^dU����Y0,�����῾M�v��?�^-��A5Pm8f4bfWY�.��	�
{�����m���P�)�hL<r�?}ϒX��ض\`�R�7��0`ݹ�t`�V�+ۢ�f����ݰ3���&�h�#~T��6�Z��$v�%���xy���	=��R�nW�_�H�7�^�;	�<^�vzM�A]��Ѕ�QUݪu|K>�{��X~�I�̒\\��74��u�IȰ����2T��L��{��2��ˣ�D�u�7Ct�������D�0i8���fI�b�ɾ�����ai����"�QK�w�r�{��*����>��:H��˞7Go���B��^Hc[F�w��v洟	~pn+�~��ͩ,(����M����S���V����UD1��T-���IA�Gh�}�*��H�o"�˞������H9Ͱϛ�;�H�4|6X7��7I��sX��K�n�����."a���+�}��*�,�e�!)}.b�0�ͼC��҉}%���p4,1&�F���;�9g�'���x��Y-���\і��<��������J�kDq�V:z��|�EK�!�q�+r�U��U�����Az�M�S؛�4�J�9X�^r�F�CG���q%�b�@�n֐�9)��˲g�eJt��˙�?�Mh��M�_�0 �pS{gd; ��jD;�ʕ�d#�o͂P��2ߜ��EƆ?�|�۪m9�k�&sz�^�些���M�ň�wa��$���f�����#M��\&Y�ڷ����"?Gl�@��QqY>$'�D�O�7u h�u��+��}�*V�0|�A��a��D0i�!<8�d�6����AhdS��p~�'dA��.�3
#D�B&�a�\*?�0�ni��P�0/��cY����0N��*����Uj;��|�������Ѽ7���Λ��έ�'|�ĩ��[*�c��l�:��"�V��ă~[�٢E[4����YI������_��0�,WQ��h!X���9��o���A��%Cv@��΃PA�鰟+��[�i03{Dt���2l����+gk�9��:� M�/v������s��o*�I�7�o�����J���� B��;�ڶ���X��I���j������ ���e����2v�UP�M�[��-Z�Ǧ��CK�`8'p�|uzx$,$������`���R�ݲ>Z�Ψ�&���M��t]�ۀ%?+m&�"Y�{ԕ��fUd�Fi�
<����1�4F��H�LB�I[Ĵ�Vq�M2�khYdǗ�U�)c�*������qz����y}���[��s�Q��B�[hh���b�A�V��M&D� %��^Z�&xƃ*��k��;�A�J>6���b��c�Ⱦi���`���KA�(k4��?dPx�>ǵ �6�`@A�8���H�q0���(B�zڨG�dqC��QGg2#vyn���X{���/t�Ĉ~�W{g�N ����]QʻL�!"q��(�A��)����W��y���j��k8
]0]Yy����٧}�x��U�!�P������W�6P��x"]��*��w
?7p?u���˙0���	��_gȲɔ\��W���8j���䉠�{��g�\PO͉9�>{�VG��V��N|&�\�⇉�(�8=���RˡE��ɠ%�c��p�A~U-4*>�Gu������ɮ4}�ۖ*���s���(��G�yGr�3<����J%))���D�U.r�U���\.]��%
��`nkI��a�N\��#�ʘNf
&�k�;�^\��������Cʆ ���FT��j|F�G���K�M�T5�,�c3,������Ч0���GO5A�Q����W��}��͂4bf��o�kܗ�5��O�M�!����m���8��K�B�é���F�֜��[��L7��F%�(�s֩.��{��������軎'*��iM�
Jr�Not}_7�& ߸�]�4�� �����$3o�������E?b����]~	��^|��V��u.h �$�[�1j�λ�E�!S*�}�a�
_-Ė���'��+��;+C �"L���jV��ؕߞ��8��=z��e	�4%���x���1f�b��0�¨v3��5�%��ènq7��D���G�C�t��ތ���o�G<�	�*�ae[*8��.�l+��O������׵��s0�A�;����������GtĠ�xM��Q� p\U}��3�����}e{�)y���o����h]#��eN�R8�32��%ԟ�D�ޘh?+!\aX�\���%�F��Jj�1��ɒ�Q�z:p��J�n9:�x�f�L��f��v��Y_�Cd�	�r������Q�:/���	Q����r�r��H����۽3�W (���
�E|}��q��!͒b�G�]S(�q/E:��X�
�����,���͕f̼��<-�7�پ������yۃ������z��dmPn�d�����ډ�#��1��͍V�'��@%;B/�@ӥ�(!���o�^�a��1�_���v��rW��-�%���-��D�D�;]ls�Dn��J���M7�d��/�U�|F��ll�Yq�U�M	Z_`�ٳ��H',�N�~���P�$~�t&d�3��jv?�	A��H��0!b
[w$�x������9�4_��ī���T�*�y�0��&*y��[�%ϱ�83��U���� ��+��A���o?��L�'b��r�|�'^�Z�h�;_����]��H�FV@W! �o�X�����J��Z�	C�F�8�J��M���5g0zW��r��:u��r�	���[~��;����v�����D�|��-��V���Pb5eW�NTVz�ζ�c�d��0�C0Tb���J�,������%��(�r7j�����,�	��[��5:��˖v��$�Q�������y�HԞ�-P�Y�2�ShFq�B���,��Δ#!縁�X��{ү*��� ��qd|U���َ�=�4�[�:�?z����E	��ս���FA��H�;�\���`3m(-��w�3AJJעMA��]ma8]'� 	���L����W�Ј|�]��l�~i�O!S-��׆����'�;,e�wY1]���E�N��V��M�,�����QCXǾj3���Ob�~����`��Z�+nM�*9F�c�?�Ϳ\ ӄ �Ea�x+q�qs4�V��9�p�)pF��VT���^����ǂ;>O����5��,�`IS�CGd'�[	����ω�Lx�d ȼ��s���'L9�,ſ�ׂ�
�ۉ+�Z�^tg5`G���r^�d�U�0���p�c�y�<`�ȣ2@0M��n�ek������/LD9�6
�wĵ$�|�I,=^A�eG0y��Mev�6��T���ܴ���\�F�
:�c�	rbZ���x���,�4���r���F�]1!�p�����B���M�B��q��gU%������%�����a���N�*mV�	��q����l8K=�=��ư�y�*C�l�)�¸q�ɼj��^?�ۈ�S\�.KXN�R�׫'EL^g8��~�:
��C8����d1�B�n���8t��-��yE�p�� Iy9��H�$�
=L�3��I�:��Q�ӽೖ��>��Y�4��
r���G��q_.��	��
i9J\>3�\�zL�l��˲��S�Q�W�U�@�8�*B�"Z_�)�L2N���
���ko1�#���󇈹��ŝ�(MSGx�Z���W쪫��k���g��5�ӜH�m7�L�����oN� tLVLtL����I�ܺʓ��~��
�m�5Gt��qC��.!�UhU�fo�E����B�-��� ���x2㍏�:2)�h�s_=��	q����a
j�15z����'�q��󌝰� ���p��u�dM��6�5n�&�?Gk��z�G"b&���>��̨�'��Q� ����I��W��Ճ�!�ca��%#ʄB����z�����,U�+��}�����v��(���ƨk�1/�$R���f�h֏�;1�ҧ�s����DH)Z0�3?�V|��OG��'/$B�7�Ѡs�͏����@g~�,֝rx!��mS,��d���M?�0N���'��;	!��R��.��(�f�x�2�1��6��g��^�Ѧ�)V�x��J���E�)VR���!�q�믢�:[D�'Dq�M��,5����~���+,G�y1E^i��ܜ:u����b����nQ�} ���x��4	h�_$��,�V��	�L���f��(�ޖ���>B*-$����C�����e�>�b��7�9�^��Ч�+\�)�띓���HR�V�fJ���F�Q�l%!2~��4�!�@UUKp��SIy�ZRk�����������h�]\b!�d8�/�@�m���H�3	�X��@h�a��6Q�|���d����9�u#n\�|D�|��Fx]�r�9�|bxQ��3ṯ}a�T��۟0 `�]��'7h�
2P�X��P	�\"�����B2��������{��׻��e��9t��V ��l�V�|���2�\<p�����N��ǣ!ld�`�t�����[�E��*��ͫb���ǉBЧ���	�j�l�����]��%�gК���r�`EQ�A��ר���]��ʑ�����._Ԝ(��HҎ�����s�S���<��&4��I~>���4��U$�9N�;j	���p��Tq�$D�O�e~��Ƴ��1����0��I^��:�%���Zw�$YQ���/���v_�ec���'��S]O4�(��W�������0�9HXF���:��I7��B����Uߨ"���8��`��$s+P5sq�ߓ�<04��	�h���R��9���pt���K-������e�K�����摯��!i[d1�� St)�"�~i����W�
vU�ļ=T-�RǱ̋J�k?U()��P+����UQkvC��;��<П�4	&��Q�9�w��Gb3}?ޞ���L��)�0� ;����X����k{���O�=)*�
��c��x�˩L
0��ą�_#0?��D����l�_8&�󲓈_�1Y���j=M;4�W�0:b���*Xnњ�}��à������2:ova�!�w� ��#']�b|�	>���wuCH�0V?�������^NUKf~޸�o�1�*^ɝ2�-VC�"������Re_g�8���ǲ�@vY
K�o�N�P���xv�@�:t?��T���(�{Q�ER�ұv�F�}L�ͅ&#��.+�vE=�^�U_��)��\��V]����+�_1Lc��R8���(��� ���6ـ�ŀ�3�mǷ���F%�c���R6�B)^n׀����R�	L�d�K�"lGӃ��E�>�H �&�q��M�4�`�SapBVjNl���:�g~6���Dr`�#��C�a%�	���<��h(��A��+����ږ�>�v�/%�"=G�Uۙoĸ��&��2�Jד8�q�J�����}<z�>��C��=��0�%m�Xţ�^�O\��{ZF�������Te���|0s]�a�l���n����[k��\�r��X���T��;�*K��`C7&����'�JF:��ub^����T[x�:!�b@�>%�#�o}xFs�b(���'C�P��.�3���Y������KB�����Z_=��ǜ1��A��OC���I`��~�b�"he�s#��8�/6�h�S�v�Q�Й��k�w�����'�(��+����x�O?0��H0�e[*{�Q�f����+Za�R��r;��տ49����
�)�Z�#ͮRyO��U��_;E��z*&oeǗ��TE�-�����hX�$��3�'-G]�ٴ�wJ-�)w�J՞\$e�p��^��T�8���-�盛�XB?A�܍�-����'�����i ��b����ue����/\�3;��Ϫ�����^c�dX���0�'��(���h$������h\Cs��^���5�h͈<����`?���2�K-���=�J��p�[ HIK�gtiqzDGl�~�_3��ש��$ۇ�
����}gNCM�3�i���3nP	0�t�����*nT�H�)q{Di�T�aX7�F�J��Oe��@��װ����N���yu�Q��˷��A3i2_��ꪐ�)�E{�M\ip�����r���O=�;�5	Vs���I��������1�KC#�n���'�֎��壠3]q�"��'JF;t8w�2ۜy�%x��-ܸc�*P��,_xVi|�S������ǂ�r��MX���Z2w
�����<Mr��!�.��~�Ż]�/�O~�DP^��W�<��t�X`@m%��hk�[��*=�z?m��#|=�[�:�8�?�Sh��!{�'�X������I��q��BXϛ�>��e�;��L�r�|����K\(�C���_ᓐ�M
�J��@\�n|�x�O�����v �"&�q-|�SZ��Xj������%�h�cB��3<x9�{/H�[�pٌ4���61cN��FR ��җ!���^`��� ��K�ߜ���UZ ��@� ��[�3-��փ؜�-���XX׹��P�X�8v>Bv9��Mc �����B@vW!�nr��9}g W�H>�"f:�[�����7�D�b�	���-$f}8	�n���}�y&�I�L�9�����5�5����zGf�ߨ�g��@���	���r�98����q�N��A�?��Ft���%+L���̓vV)`�>~�������ѣ���^{( J@�B���w$9a!L�-]9&�2�ߋI��p����H��=	l�U�,���W��ť��6?�,����10�#_N�D�ACI�<�?�tzy�{����BY�r��WT��Y�.	\Ϥ(��C�@����	i�ң�>���2u*��[~��0[1U���G��Yt޹,ڒ��'3��&�]ḟ���>ڳ��uXs_�Bف�in����dr66<��	�ֺgU&����Ea%÷̂5y���8�l�R��g ��R�J�� �^?�f�paCŢ�\Р��*����a��qi�'a9���z� s+í������o�۴مiZ���Cn.�k&��<;�ORQ�X���$]�c����ھ��9����n͜�=���'=�vG�~��Q�g�������)����E닍�Blݘ*��x]}H���ٝkt(��H|w�*�c޽!ȥ3`����d�@'��p��TX�P�H����	�~5t,n���N��}���X�8H,�� �q;���e��be�֣I�0��F��IP���W�`�@AU�Y��h�7j�AZiՁW�[�4�R�{����bC��V����$"�]8*W�B�1�b8\$�e�Ko-u�;���O�\�~�\�W�vfZi���H�	�/p��gE�Ь�J1��u�v����aЈ�*x�pF�%Tv~m处��z�������)�{4��e+	2xs�/����Uy�)�R8
����z��̳��ߔ��4~
���d2��sBH�C�(�++l�.s
�$.��%:�F�s��ؘ�%���Q3����cf�d/GP��n�?�LK������4�Wr�*f������7p�c���1�;\��_���+u#e�VV���<��s����92����|�r6�(���h�H�gڹ���
����_�v�Z�2��/��u�&���"��<�q��������h��y����F{�3v�(8@H��KFL�}sJ
��;t$�'�	��K3:�
;r���UjK2�f��^�����y�&�E?{K����߹��z�b�'a>4f�~Po��jQ�(MnP���i� �b�1�ō��_c�s���:�b�A��Z��H��� ?5*J�i������Z��B�qp�WS�?�6G�>Y��?�)ZK��2�ZЄ\��QVW�U����D{�+O'��SmW�6���+l��Ӫ�e�q�ك^���>�楅sY�2�js�0%V-U��F��
�(W�J?���1t6��kbߺ���u���5~�XP����(�e��C�=��T�Fda��O�-=~Ƿ ?-]iC��t?�[��{HԒ��9�^�
�^��h�ĕ�ۺ�m��>�P���ܮ���~�`$\�������5���m�!��~�Xg��q���TbdK^�@Vc��-�Wl�z�W@�Kr��ڒ|V��H��gM�]��z_��f;]����f�8kU ��e|��y��o�2|�-������ߖ�Yr��#�W|,�=�rC�Q"�琘]Ο�#��O��r?RpɺB
k���l��ƞN5���5^�bDӱ�O�ؠ�H�i|s��򠝉}~L�x�7�3$0�X��b��~~并�[�ƶ����&I�<��!'�����O��N��*�xy4��IlZ��̌u[?��Z?��o�~�hz�N���5#QT,P�v�sh�uM���8�
#��b)��[7�L����w�$I��������+�U�;�BX�����Q`�	�/�6EB���#S�Y��})e�8[GO:SM�ѡ����X��nQ�pA3jH��{�%��J �eX(��S�{�b��q�kP��|	K���ƥ����tf9����?��t�hg�n��Tt.��.�Ssv�R����f��=gh�2�ne�:E�IJ�hL�% �����P�����vT�|hLL�D��5��ka!�W�j���ճ�)���A��u��c�6��EU��q3c "���m��t�f	���0([w�.���f�5D.x%{����%g�0������tN����3��B�Q���W⌒�@�Mj&չƙ�f�gs��6l\��FyMJ��{"-NS�E}���#�pX$Tp��"^�}�?���'#�$��6x��B�U� ���ډ��%wT����$��XU��G�)�b��.!�����<��?���ʼ��n��S����;T�,���L����2~�u�'���1ʄK��zKd��ͤ}��KU�s@�*}�	lץr^�҆���] ϰ-ड़�2������ZL����nG����V�ǡ�V�����	}Sp6��S����"��'b$�p7P� ɝ�Q����oGj�p8�eI�:�s�B:�(��v��E,^-{�1�
��~h��0S����?Mb�N�K���[����K�n.����1D5�oex��+���~`��D1 �K��q�"�����c)F'
��)�>�Q����C��e�W�F%B�=7�V�)���8K���K�;�#�3� ��� �e`7���޾�'L*"�*�n+Aּ��<j�0��UQ�#�e�} ���xR0�l�jn\j)�-�����c��V:X�����pwv����:䆪��9Չ1�dZcm"͔�3�DtG��isUV�A<-��Bfn8�V��l���P���]�euC�"��ƙ�p���&H�eH�Ln�Ks���Q�1�l�I�tڄ'pB�l����Xn�&4�5�P�054�t�}W�-״l�XF�6D�S�����3��:����G}�ҙH��g�D7ʑ�
�����^\�cz�4aBLp�::�lA:�����cs�4ん�M�I]�}�t~�~ݺχV��C��'Qm����j�"#K.у��A�-?q��ݣJe�3k�ƺ� ["K+>H�-Օ� ��>���S�K�e�i���*����n)#Eѵ��v�UK �k�E�Q���v�鋅�H�,%:�����sGWYn�] ~M`��ڲ�F�)j_�U=�!k7��Z#�Ef�:����UK]pʝ���:P�"����4��o���4�?y+�5
���Q�C��-���.�B�e]6���~�YU���v�e����3|�� ���c�U�k�~���pj��\���'Pѕ8���N�"=3�~�������mt^��PL@v��s	/�3ff-�i&��|~�k�
����v�_��J�������l�,~�M�a�b�6�� �����O �kbt4[L�]Z���=��B����teR���38+(:�����D��?ĸ��o̖1�� >jw�d��3ƻB.�'c�X�E����O|W�*�?�T��)����^U���|6�d+]�K�Y�AB��󤍇�I��|�# O�,F���3�y�����f�J��:�����m������\�C�yC��JHv���Ɍ3����o9D���~�x�ѝ#�L�p�VHj}Q���<�Ȱ�R�}��@L���o6e���*]��x����B�K(Qַ��H���L���s�
������y=%8� j|3}|�x������Qh�G �p5E[��l�a��"�WU��v�@���˧�P5�ˑ+u��_�F�ĪG��l?̳y���sT�I�Xh�c�GM�$�%��5����9�>�ؑ�HpҐ\���j;r�J�
���B�s����G?`�IkY�KmA�
�f�V�U�F?z�B��9#�m�����s���pP��n�]��f��d*m�.*�����S��N�26��.�5QR������ ��C���1s�4�y
�0�R��Y�3@Y�!��B[a�/u�K�b���UL�93P]�M����O�Z�n+��0n�=Q�-���l0�L���s;�g9$�<&�	�|�Ǹ~{+���p�Tsui�+�~$ItjTj�{_<�X�Y#!	p��፫�J�̘u�s!K��n⑵���Q��[�P�Xo�츄�G��Q�����\ڡ� ��m<���]�^s��Z��.Y�7#ۜ#=��@����^�DD�1Di�]�9��Z휰)rU�Cӂ��a�arwm8v��H/��g i�q���R����N�ljp� �`0�ºn��	��5��lִ@� <�ʲ���{O�I�\���r�>;��bO��2�gj�{U�Zjo�/[r����"m��	����`�� �L�ny
�E��Rw0��I�����*��z�fd����X�����nd�J����=�≠�`|��t�A�&o�daf�Ts�%܊q&���M���ߚ1�ti������3�W�L�^#Dl)��B�.es6`�
e	'�����W�mϳ�e�ԣ���k��%��P��eȾlo�ض>r��2}qb�Q�˻��뮟� qd��#n4I�T<���i�5õ�IS��&�c�U�P �ͭ��h�C1]9ʄ�J�T���kn�qq<�%�8�WVg)�p
V�)���Ӄ����l�R�yk!ʸ�=8Y��(���$���&Y�;p�v�� Џ?�.iT_H�D�x���/B�X9�pv�L0��)ׯL��^?����y�T}(�N�G]��B~�fЬ��~Ĕ��ҏ�5z��ᑟ�/�nlW���(��J���b����F�����K�A����<K��G�q�-jE6�O�j�����ʫ<*��cUE��5T�`�h"�gi����~�>rఴ��
a8A{����A�����6��3q�%R�O�^�\�u�K��#��n�u7f���ɫ�Et�ç�N�c��ٷ�#z�U�rif0K��F_��!��6xǣ೾�)>t���G�Rŕ=�|#��k"Λ������&6h�'LZ�NS]� �H�e:d��������14�;��}4"�:+����Z�OV��}��5ތV�i���:�t��9�����usch��l`��;�.e���u�Qrc
�m�M�pL�� ���IS��*�:s,�p�]Cp�zV�j�M9�'!�hz�T��o�3˶<C���x�	���+Yd�n���<(nM���0���௡h�P�i�%�!���2����X���b���g�'�Q����uǅl��3t��՗x/+�$����W��$"��(`���O����u���\'�3l��`�j]$l,��v^B9C�����B�牒jZR���+���� R��#*CG��"�
|�Nh��\�]I�P�ސ��2|�"�9�
q���xh��kg�?��{p�����e��������>�.߹����f���6/���Z`�}��*ձ
�)�H@My­��삱��[%�+����]P�ڀ�T��=��qG��MI��71��q5�����J�
ƀ��th;���y�s�N�o���>A� ���E$���1�&=�ؔ�7a��t�,�*R;`��
Č3~C��z<a��;�hH�&HI�G����}��������.���=��G	
��Y�K�IF�nǣ%.�<ǩ@I�d�nB-��W��9�4����pF�=5Z�;Adg�ت��Ô��|3[�(�L���D<K!/��)�ޠ�.$���{[�ٱ�Y1#.��1h4��W"9�-��i���<��vAg@i��@3�\}E�����h��8��!�[�W\S~G�P=�> :R�̠��q��f�t���]#�)�����}E�\��N`TR��	H��}SQ:2rG��)�[ p��iu�39/^}�e):9C��>�>�r6X���٠�
{`�'���5=�큶���:8d(�V�Q�^�������a��!/�f��S���mh��9'�Ø��;-??˒��Vx��S̗/*D߶�Lyi�G�Te��K�̿xKx�ZOF�6�8ǭwV��/��|�_�RGq&�ei��C}���]�������U��qA�^`g���}c��CX�"�&ޡ�T�Tk�W����"(F?�46��>�`�h'�i�7��B�<*/�0V{i��0t0TjI����QSs4�-��*�,�r<��	z�6��tj �s�Z��Q�e��[�E�D-���>�d�w�%e<b�:f>��$�n�����i#F����͡`E�7��`�+��`b�e>G�P�s��7}.ǬH㞨<�R�����"~qY_=�&A&XK�����j��	T���L�q���jn�}?
#v ِA�z��r���*�K��k9)?�y��޺|�f�ٔk�Ƨ���uo��B8���)�wK�8[9KZMJ��j�Ƭs�g9��o�}�3���&����)��O�vC=�x�c@���6��#S.;b��ݰ����vu����t��U��Yժ�.ܚ@:_�n�(�NP���=ZG�"�vMqs+He���7�e�K�;�	5Y�n�c��,�<��TT0�ʢ�B�/q���*D�%���Vp;��:��5ro�4���.�M(�7������@;>}N=�i��<kbh��ܲ�*A��(ݯH�����Ge3���o٫~f��5.��c��YL�[��Y�A��Q1�1L��^����ghzj�����>b���5��ߖ�%��7:�?e�B瑟bu�`2�ls���w^�+Q�<���&�j(��ѻ��.O���ө8pׄ�0
@����*3~B�&1��]����9�:,��N�a!�i����I����4�1�������4��Z���u��kY]�4��5�O��n��&:�y������g�� �i��:�2٠���6�ӋF��.�P�xG�Y���EO��:��TC�a�3��vbyL�������#�D�31"�)6�j�/eI�)��K�����������ӚW�S���T��-.�Z<��:*�>W�^������s>nP��Y�i䊼]�y�sE��� )�9Z&���7u�6p�g5����S0k=��ᣤv�I�Y����������e�5Lt�\�����V�Z[f+�u~6������)��4�v���?Q�	܄L�jZ�~d:�V5��5�|�8��T�Oe��iK��������s��t�-i��T:c�u�25 �1��!��.�b�X�I�*�̡� ��f��[3��(R��=A������y���b_���� �4�W?Ag!��{l1Z�eq툎yR䔶�9�)M�3f�B)�V���>F�C�Z�*���>m����jg��rR��ƜqS�.!�X�S�������Q�"��"V��J�(������>"�"y)0��V-��v�#J�8Ch,�1��=����M��x����_�,*E��P�R�����q�~ECT�x�ˁ֋UҔb"�����V�ǳ�bنv�$C�%�AڶN�X+�7>����/3k$q#��;�J��&6�RA�F�k�B�����Q��Ī�1[�N���1z-��J�%j��j�a4h)k?Ӳ���f�K�A�8�'(MCX��rlF\�x��7��RM�`W�)EV���*觗�9��g�㦕���'f�ꦺF֚q��~d�6��ǌ�>�7���qW���U1@�S#?�p�4UxJKM.q�/
�u��C�oU�%(�fD��Y (������Ǩ�~۟�4�>��s�]{+�
�Ȏ9�%����p���E;����K%]f�RA�>Ą��g��n^�����Q�@���*P����q&�P��'e�n;�4�vy�2������d\���XƯ����i�HԘ�����Ǩ� �G.��Hu�
@�8-v�8k˓a<
giA#L��_g1\��2��DjЃ�V��Gb����9��� �tG�j0�a�|�'�YoW��O�!=�=8��mbWB$�j�[��RԮ��HP8�����0���w��z��2):� A8��K�K��������ך��(?!w�Mh6��d��6�Ew��j���p�"(��	/�Y�kpp�~�d�'鱥-�M�U��d�.${�P�>�dS-6���8r�"a��ZO�?(R��k�0@�����Q+�l(�<-���{�R3�2d0�5f��b*i"GG>3*�ݓ,�~=Yc݅�Gw���y�N�^���kpE�j=����fN��ެ�\%oy#��*w���p6tcG��W�i��G5�z�P2N|T�*���\.�%@k2z�!���a�`.����V�LHqe�~kn���_�S�����v��(:m'�۲	��˖�"����*��{&*������wa�>�,���s��pҗ}�BA�hY���$�m���X�3���7e(���Sx��=z���d	m]Rז��aD,++��].���ȳ_DN���a)O-�"%Jףrg�t��˹�C��9g�`��U%�b+;�r?�JIVL��4[���,��O��*��h��pԔ���_i�f��D�J��iE����NHd�t�-\�=�j�il�04u�)煶��h�<m��U+��IJG�M���x����������3�y6c����PNf`,kMYN�dTM��<:˫�^˪K#酃�����I|93�}O^���
FaV��v��)�E�.�;L���,ײk��v���]O-R+����oS��Q]7z@)�3}�U^�C_3�h�G���I�� �랤�6ل>�fi^�n��I>&��$�ެ�olm���:��0̸��\Z�w�	"�:�Q���1��^&kr�G��ݪ	�LF|B�n��f��-.���ؼV��u)�IH���\]s�#R�4,��4PG��߻���N��@�O�IM
���V���Le
���wj�u����3��:��� ?4��e��ۘ�;���Q�xm����Grc/,j%8�7G�#�8�M�.d��A���,��K7(M5�|(/#k8MM ���(�-��r'�)[)�2�#I�ȸ_����×�"`�N߯p���Q�7�g-���YF�ݚ��6+�d�
L\�����o��c���М��S�����7�+i�����\+���#��E�l���S5�O��#o�rYG��ۑT���8�Z-#@1�Oy{�'���O�['jb�J;b�`�0������hr����1Z Ǫ�Z�@e���m����\ϓ�,��g�U��XQH�A8N-tښ���#�y\�N����/����Gw�OK˕.�Pt?�W%�L�,���0T�.k;)�B�ʋ��W;H����3�Y0]
/{o����K���A��ʙ����P�9]?l�,�{��4�Ja�C���G	ML��h�b�p�����{�^6+Y1��Š�������k'��==�F��T�@��Q!^��럑>�!^2UO%��H3�ζ'�����U�&n�d�B��>l(+�*�w�ʠ�vG8U�� ���U?�3��F�����Q�CvE}�� �Cm`܇L��P��Ӟ^�8�Aߕ��Rg8A��?�]�}�|K��"�gU�VMV�7�_E���[_g
�XF'�u�\5�;�	�}��-f�:q�� �/Ԣ���r��(/̓#a�X[l �?�_b�r���u�],
��]V�@�����򃪻c��f��Ӣh|t��v��G�-����Z���;C�XĢ�������ȝ�;��ƭX<0HJ�<�|'��ĩ�W�frC杤�a�$�t��jа�QsΙ�N�1�k�=�,ub�P&zu���%��Eo��`LLL=/�
��[*��e3ֽlH�^�v�i�D-��J1��q��KѤI��}CV��7T0��u*�>����Ǆ{dm�v��ا�O�#*�ֳޤ���w�8�`\�y�I�gჴ��dp/t��3Wm�*8�2h�-��@�,D�1����:�)���	<�egS�11�m��9��%��]ᲃguR8��Ix��id鬈o��r@@�l�u9�dr���(���r�QӰ(!R������'�w��i}�n�R�8+7i�B�3^�X ��(�Ϥ��~��L���wfd{y&�[U2��R82�V4k{a&�m��̈	�[=�j �sg��%�9�̨���P�3	rl��&Kg�Ԧ ��W�b8` �p{�$�^yp�n"I$r����p��f�� �H�4W����\3��H5�u, �%�!�P�N?2E���v���/I*������3~�)^�R�@�=*����{p-��M9ޜ�݌-�~�۹Ӽ�>[�.&�i� �J��Sׂ��7bf�oH2��cs�-�[��� 9h�q�ġ0��KP��+Ljw_�E*խs3w�U���B�
��>��J��)�����c�(��� ���鞞���{�9.��0�>d7D������םY��rLY�}�I�I�
ƕ�7,�ߑo{���ɿ
�i�/�W#���﹉����J	4iC�4X/�!!�h��b*4;m�s��k��h/Hޕ�3j֋Oi��[��^��'���Ɛ[_�_z'�u7ˆWU��T��&�7.��P谼��'%��v����Iw�p@��3��oħ�jښ^�M죸0ݙJ=}ֹGء��J��ӈud@��^%��� Рx\�k�S�H�o��Y�5�ƀ+`��=S��z�Z��ğ<�!!i�W��̄�4X�:z�3����Tw������rJ��j�ڹ���2���ɏ�C�ӷP��?Ui4�34��?��Qh1yz�x�}�ڃ����/59O����v��ټ�A<�<�i��5Vy����6�D"2�D�l�3�3��#�E�t,&=��4 WY&��ŉ�5|���M��K"X��<H�i���:ҸjoGO/��Ѻ���Ά'�4���c��'�����z�V\��
�n�2�$Jn_��OIV���uUJ�kHF�i8�iTrC�5}���P���:��Jl^r�����&��6�R:��_]`T�/!P�� b��d׏��z��=���}r��}�A��t#h�Z�FK�{/�_���gOu�/�m�4�
��l�����a��V����ʭ��*�X���7��w��@GŢC���ʆ��"e)��� �R���s�v�1yP����	�"<����=�z偫��\�>����i&pW*����Q�'x�.iv�L�iI�F?&���b�m�p_�E�'��N�a������
�F���垅<��x�O8�&�ǃ1��l/̡4����5g��j�:��g��J�*F�H#~Xf��R�]z���$�t���܀��`��;��i�$�A(f�*S>��R��*����q��:_��� ����%P��9�������R$sp��٦��߮�)s�e�h)��V��X<��CQ�]�����^�Z��|��K�'Eϲ�lC�ڪ�q�0X�cIQoj��~[�DV0D��#Do��|�B�?��8G�E������3����K�/uSh39��wA�	{̦��}X���*L���b���Z�,�J(?'?����sn�M6���@���H�^���P���{�B�å�| ���� 6���A��� }I��T�4��#$�m6T���Y��'G�~f�&Yu �LdI�C�b���:cfϔ}����rA���C�s�TE-������Ssڣ�FgzS��}�S����{M �>�S�k$�k ?�����N��؂�]�N+@��)@��P.!J�=��:*d���������!��nĥ��u$M���H���I�°n�HE�c�������QQ�y�-�=�a/���,a��ֽi�� ��LOE��U���}����K�e�#����~?�@�nB�wV���;-ZsQHj2}XYcT�=�l呛d��	�t�dHl3�V[�Qˮ���+K��`��j4���M}#���ݎ&�A��ɈQ
7�@�������	���S!³�4i��f���F�?w=�<4�?�������������=L��+$�|��=��Foif�^T�,B�^�V��u�����x�O�� ���4����J�����.�4�3dr�M��#5��GycQ7��y��Lac��^fj."����v��li��8W},���|���y�|�kZBVo����\?�` �4���B����Ⴟ���ގL8��gĜ�`c(�i���/�A��Q����ZJuߵ����S�`5�+RܦV��9�$1���!:bh�x�N���q8����Y ��^�LHB �{	�`���6_k/rN%)���${]�j��<�҄!�;�\&S�k�������	؅��++8Ł��ZG&񜜋�s(�v%P�k`�����+�2:S�4���'n9Q�ֱ;�oY��/�|E�z'�y��F���!��bRA��Oi\�?ЭcV��5����eN_�?|꓀	2�����M�"I���g'֥���|�K�_SI�"�D�Z�u�ӏ��\U����}f��P��1��
v���/,�=>����+�-�=9�7Dl�����{x�+82�_ç·��E�2��ץv�=�O���^yGz����0��6����嫀����H�J��HC�Ń������^� �g� ��Y% GaA/���D��Xٓ6A�Ж_ 9X��d+g$L''������B���_<�.k�Y$:�גl� :l���1��g�i��{��~?�,��e���L�.�`�V(�Q�M�:�r���:��n#$����p0&�e� �=�}��CP<�h�H}�=cO�U��>T��h�Jle�%�`��-��ˆ�p1��G^QD�z;��&˹��;�%�:^?���ǩ��^12�Ǖ+���8V��)F�@�VP�'NhJ��ݺM��^�7\A�uE�>t�8�=|y0O�b_'mqU�k߸pH;Gdxet�L��{�T�"R�������}�BY�׃���PO�/�����a����:������G�)�@e�@$D�J�9�����O�Z/P�xĳnQ����kRct�n�݂i��,b]��ݺ� >��6Z����!��,b6�5!�$&t}|D5U�m�Cץe����VM�W����x٫V�2_߮0�,��"�+K�D�Y�� D�h�g{n1�D@R�QC%/�A�F����rw��a-�k�ܧ�P��B����_�j]�c�%U�W�֎Rr���1��}�3g��ƃC(��̺coꅟ帞-���Z�`������Bj^�!=�N/��!MƩ��޶������h������2I�Tj����!0�o��ՂXa��,�F��6�7ѡ�˒�q��㑝C�/�����Z]�rv0��J~ٚO$���''{�^p�;l�%Ln�"�sq��8�Hr��}�� �3��?$\jLL�JP*��{VQ��k�FZ-�`���z�A�c�8�9'!���7v0��rPze��w��}���0Y�SG�r;��Q*�`A���h0[m�XB,��|'JaE�+@�R�n��-k�ee�DY]Z�W�X�Q��t��􏪆����^46T�Ӄ��Q]�AL����B��vd�qeQ+��^&��y�7a{
��+1�C�s�;�j�/&oÆ2�����{�,f�О��R�{�-�My�h��`�����:@�*��%`�;���<�?�!q�gc
i��l\�����pY�ٺ���d+p���)�J�e��J�#�Eye���۰rd��2�$[A-��'�>sϸe�=��D���v�{Q�>Ĺ�@)�����56Zΰ��ʞ{B�t�ѱ)`��`����[N5Cip�����:��A��i���C�3��H���x������G���!,r'�v�#հfd7�B*�{�Б���9w��s�|���-g��X�]�zx��0lߒ^4[
�+%t,#7�  70�@�t�������զ���|Yjz�Xɮc�
��^S�7�7�^�o��Qf@笳�K"��,�%���w�$��N�jm����e�&F��[�!pCU���5k�nd��c����[kt6��P����$v�X?�ut�6ܿ[v�$�7> ��`��,�(qԅѻfS�A5����`H�;,����V/,88�?�s|(��K"���1�mu��F��� W��v�v@{��m� Xo(��cx��%���5Eob7���R�bbP@�k�eޕg��@��H���E� �F���9��s`6��Uu���ؤ�4���ϋr���z��S�h������ �����H=����j�S�2��~�7�>�R�&.�[c�w�$Zebt6M��#< U�����+��o�6���[�DM>|H��;���	��������}!�>�!��R�m��&��8���O5*1�W>��h�t�#F�����Ic�A`Ϊˎ�:G�n�9���[yy/��ڣ���r{��礴�\�~����0�B���*���x���SG9^�*h�z?#?�w� 9g0�oL��@��y�^`ॸ[w��$`�����<z�c�@�?L�q�GǛa��iO&��M�]l�a���(`�N���e<`��
�7�>_�j�X1/#W�!��Y����lf�N��# o�~�tt��WZ뾕+5��g��[�b�[�h�
�b{M�Щ��l�bI�^����s�E	H�GE�QF!����A ��y��� �:� ��F�%P�J��w.���i}|i����1W�@��_�ĕ�C��!e�6����$�xH����./��r�9>y�G愅sE$*��툭�s�N��G	�a��Qv�9��8�j���T��i��Q�4I'�6�1�{��F��i������[�MF���iܣU���#�%,T��Z��2g�ڍuY�Nt#�ʷ�!�mP��.�ʉ����R ��$���/����@�����1�`^:Ct���dP���Ҭ����@C��ac��sS�p^d�ؕV}�TZU=�,�"�E�P��I��&'ܜ�%�����5�ǈ�&[�z�(���v:�Q����֣����p���D�d�<D��"�5a��4�p�K�28�cm��S�{���Б"/�NF��g1h#�"�@�JV�-AT��#�%^�Uc���e��Q]ƀ����YABhĞ�K ?{g�T����T�֨�r�
fP�D/�n�@XvY�E�{e6x�kj���X���w�m�t����܆��Z�4��y�Ba�fu]
X�`a�X'�V������Z������-9 �S@�]����5�s��@�����C�n�7�H�lZ�OX'7�|$h�f&V}ԑ"�چ.��ޠ[X�N��,���w1N6��c;���o�G\�� �����t���>Z��W5r�YiI0k��eXh�Q�
���nb`7�nG�ף�6�׍,JH�� m:�Ϲ��IR�	�t���<n~�b}[yB�4S�o���N�5�I#�.d	�������63�EΙUʙ_o,�ZB��PGc�t���#I�k������{n@�f9��:��?Jy����P���^q��:�5�����\�)1i5�|;���0b$�z4�`%��WQc㿈���{��?�2��T��z���̡���I��?�:��3�W|ȼ� r�mA���K�x�JH!�+j	eh����T"Ý<�j̴Ġ�S'@\��R�/Վ �tb��|��_��c��t�>�NՋ��sBfdɅM5�"k�x��_�й��N9
O��4}��Y#�P0�p�|��L���R�H��Z%5<�Ѯ�+�6-�uI�lpN��y�rꤠ��A��4r�?[9��Sg�� �ù�'A*�c�@��yQG ��e�s�k~D{�X5g��*&�hn%m+nzi|���{q�����|<���(�ޚ.���A5�Z�u�R�,�x�)i��L��mȰ� ��I���zr�������F�+�>^�����ƥ_�;@.´�zk	GoN�g�w
4��]΂�hn��� �c�:D�
[*���0O2��r��]|�̱\���Ƥ���8����0uo�XZ-ۥ?~�r�"����s*�k���gFhm�L���s���1�Ï��3�Uh ��G�-�;ut�%�m���S�.�t�k�>)?��[�R;�k�v���Ʀ�/Lld4���MUDZ�B"��OVU���[�'�5�����?EJ�]�Ϛ�|��8�Ր1SW~p�}�U�=��Uu*��L�6Md���P����F0�&J�ٔ�d_3)uy}���m%�/8��j��7�_�)	���Q��Өy��$��T��
�/�(s����ɏ���#��]Z�`�w�(_�p��Yp*�Ǧ/�+q���/�;��{g!J �GH���T������93�(�>����с�ڮ����~�{q;Hl�O��8���N|_��bO�����O�#8 Ď�;N���R�z�� ���iN��[�.�!��	o��K�����z�3Vm��N��;ըv�Z��a@h��"�X��IK�M���R�ӡ�_j�D��jm �<ڋ�Ó�6ì�
6�y	��"�.� �Ң4����Z։$�f�>%�r������w�L/fW,�M1\5я.���Cg�>�pT�p��`KI<�uZ��q�	*ڢv�<:�l҅��k��X���A��M{ig�!P�:B��.�������ִ!�8L��l:~��ւ��z�Be�;�4Ro�����8�=�b͖��R��t�<$z�%*W\o�&cF����p��a���(�I���3̗�/9�^�fbp��DToJE��������S3:dO����7lۮ���=vJ�P)L��	$����	}A:�}n{�e//�4�8���V�i��0Y$�MX)�����ֱȝ:�*�O篚 #0k��%a������������!nQ�b��j���.����)���9e`W�Yl9CN<�%#7?����[�ݟ=~�D9�CcZ�%�������zA�Ɠ���*�H������.���T>FAN���@,b��ܜ�6�O}}w���� ��Y?ì3��,`<�+�G9�+�Ԓ��f$�S��汅p��S�Z�L�A�ɼ�M����g��g�E�*ʾ�ó�1CE3@gdP5:����<ڰN-�v��d)��W]o64quf�eO~���y~"�x�Q����T�f��AE�<]	j�X.�w��׈^Z��S��0���o�@9s�W����j�i���ld�_~��bw+5�W���b�戩�-Hmr�d*x	��J�E?�I]ٿԼ���`�n�ק�I@�-�~����Z6����ߌ]��4��r�!����K�γla�c�㎟pd����*���/Dێ�ֹ,��?J�{����1�l�P�T�^��`��i'�����Y�� qn���b�,�o'�p!6��~Kr1ۺ���k
8�|�c�RY�߫�0�G����<��O�p�!ӣ@1�AOQ,:��;U�-���� �qGi��v�j�w���Z��O쨒wL�y\���d���x��Ӂ��3���ߦ�|K=��'�4D��Gw]bQ�ZQ1�Ksf��5����T������v�V�'����B
7c�_S���|��ժ�X�3�'�B��q!w�)%`�i�Sh,J�&�tǋ�[��{��-(�֟�JPVze��>�S��s����0��v�1�ƭ��7/Yc8-H�ʴ�;&`E�0?O\=�����y�3w/u��e��ȕI:Nr�Ϩ.��o@�fȱ3�ZQ���s�Ԧ�� oh/'`��W��ݵ��os��4��m0���L�0 xW�����D�H^�~����Yeϸ�1f�sF����]�����V4�Y���5�£��JtY=�yM�$Q�#��¶;d�`�c�(c^i"eTg�<��5(<��:���*B��S����S�U׉
�,���m��r'���ѵq�گT)���Cfʬ��N��z�B=�t�͇��-��ki�\�h�Ul�������M�/����_��i>�D�b3^]�~����tv�5����m'�ޟ��D �Z���ӱ�ס\�7�n�����&Ųh�\�$!���p(B�M-T�w�l_j��O4����A��������{騬\�UNe��B��݁�ZN#��9ފ��R���j��0ý.�]�w7��Ų�g�`f5@��	5�> �]��m:�|$
���mYȵb�l:Ow�������ΗC�&������ܥ�O�}_���o�ˣ����O����L��i��s�2~��M �2�[I
�B	���B@#�;ǾG��&Q֣V���.�����}^��GԠ`8:��Ɲ������ׂn�y_��kU�&|�2��Acr��iI�<HS���5�*��腈U�%5S�qn�["�9P"��/�X�J�TT�{����H��;6˨=E�(�B������	�b��M��!`�����D^R^�����y��UD�|�I��T�s8e��$��H� ��+�@�Tg�H��~�	Ў�=T�-�s����#��)ku���PdeY���΍ j�ypT�e+�;P�/$c:���EX<�}0ݗ�����s��C^�eX��6���c��w���"��XE !b]Q1m�G0Әv6L��²�p9������F]!�_5�v���<���xhVww71�[8B	�X�ZfG�xx<:�Dp_>FV������.w&����W"��Uos�����|�*�o��G�1u.�VsJ��^e\`�ֺ�^�M�W#��_��YG�s�]J�*��fZ���Qۚib�v$z%+_x!hT�Tr�c� ��J�η�&�HI�i,�R��*]*�2+Z�t#�����������E�,�1�'��8'Z�&5:W��/	�Y�g1�f���k1��j~��n�.<�>�G�Vٛ����G���;+�C���T')��2{����
�](�a	,ZA!kea�k��[��Q�m_]��⢵�)���M�������L�P,�n���;��<=��X���}���^�զ�y��F쵱;�����k7�	I�o�p0��&���6h�0��L)�eszSN�D���j=�d����t2ʇ��ҹ=��k�6�e(����l��:��Y����M�\�]�3_m�&��mB��4;��V����^�:�9�Wd�0~�x�>l�h�F����2v�U�ah��{�畺�ܼ��6�Q���s��0��Fq���q۫X��{}4��n��p�v_�tE���-*Iv�Uj��x��?�Ϡ�zI ���V;��D��܉�<�5�c��e:/�T��Xώ�}6�u�EcJ�:f��.�3tI�%�m�3n�D-�Sm��q*��<�a�U
C\b�� ���e�q�1΂�APM����ǲ(��t�3F���G��`�=�� [�q�7�^ם ��L�M4�́�HM+�ୃj:�'�F%]��t	����� ���9���G�'m�:�~��qsC'�I�����> ���$&�y��4�,����L�����R:� �xV�3����]���R�X{!X6��SM~cg世p��7���w<�o'�3��s�-�?���o�\�7�t}`98ž���O���:��)�G�j�a4�����#��#����U3�M�-�	�"��p�D&�`�=���t]+�ƶ�o����)����%�����Gte_���T������oB��-�A����1A�u�OW�����$E�ʼ�l�ᩅ��]�5KUS���G�k���c�&�������%�$�g���H��>���	��S��q� Y2�!��O2�W7v���[Kv�zQI���4EKS��ީ��Zׂ�1������Hj;�]�[��Fy��X��9'��Wsͷ�ٔ�k�`���k2��7���ny��6�\*(�Uu@2��m����U�e^�Y�c��k2��{a�R��vϔT�Fs�$	n�ō\R�7��`E]�N�`�.?�b;�����_0�)�.Ù�3u�H����ä���ِ������׌����Z�C�H��Q��s�a�9����<ؒ�4;F��T�ɫ^�E�QS��
-� ��7߉���bS2�>���o�p�T���=� �̵��oQ^�eY�@| W�h��?���!B���d�B������e~s?X%p��>�B�k�wb���1�^��}�}8�{`I�ǴC��L�����ƈ	W��V���샐�̹PeQ���{D���UH��?�X*�/������_��w?��3�Ru�^	<ki�ZF���>`��6
��v����d��!��֕0�[�ux��#xM~-,�l�Κ8����������ba[�ҐO(�6���p��RM���`��]j��Q5�	=K���
�O/�,��^I�`���ۘ�$���se5�Ib��p��@�@����߀����v,�iA�|^�p]���{���,�h���9��iA�ս�'�V��	�v݋����$��Ȩ���⥉��CT\*XuO��!�Yq׺��EZS=�D�v~������ʮO�@�C�̔��0�6��W��^l fW;l���� ��iG�����]��u[��K�FS����ړ|�����VWQ�<o�t���4r�L����
H�Mh28��~��,6���3_����KF�yJ��@31�}�:�����R�X)���E�Z[5|��~߈e�9!��sl��JVA���D�ڿ�t�P�fuC��X�TI@��|l��4}��%	@��&hnU@��בY�*I bʅc� ����U�O$�g�Nm�S�k�W�W�kC.nXv|��lȕ{��� ��(T*O���(|� ���|���ޢ���қkr���)`=�n�7����abl��ø�u���}���r�7�uR���u��΋ϯBF5B�\]��Y��}3"ߩ>x{�B�p�Jy`g��	LWN����'�������8�l�{9h�4p�F��w��1OaW�C~��!r���h7�]��&+/��*���x����YǭW9is:��z�(��FTp�h	���{QG-т����� [+q�s.�d���]��[{����u��9
o�� 4Z�&�Ţ��r�o�K�)�;ۓ1�U�_�^c*�.9yom[�0>)�%��m�DG��᳡�vf�G%:��7�����a�\�T,Ĕ�3��o��щ	����m����/	)C�f�e��QHՔ"�VZ��阯� &��Ͷɞ�)���W�6�v����ְf�[쨢ᦀ�T�HC�q�{i����l��c���WM����8bGD�o�@�3].�/�(U���D���� ��f>�.����|g^W=X(Նk���^�{��I79R:��kV�WϿB���,��R)��������D�4\j��;��#'�����Ԗ�j��إ�ګ�V�Q��a���t�OPO�_���Z�m��S�^+��랳��!�����L�v��ψ`���a'	��5,�d���:���R���7�j$�V6K4A�T$y����@���$ۭd�@��Ĳ6g��sZǠ�<�6���b��Ҵ�Q�[r[��SL Tv}���]�@s5�.��?����M���`�=�R����±�rO*-c��{W-��Ej�����eG�E�����h�A�PJ`8����F��Og�_��vxO�[ �d�2���G�/�e���\h%n���6�;GD �q M��-GM�Y�2qbn xrR�{�����U��g^�m������r���4V��>���-�+�����(��0��T������H�r��J�KOݺ8z��kQy���݊i��J��8w;fd��G���� ��sČ(T��ReW}UѴK�Ju�C	>o�a�3C{��W��!��7X�Y�yÝs,>F���Db��6(h�/c��9cҚ�p¨6���o�#G��D�W����i��ѧ��|>9�n�D=m�"��}�����r"�/�m��� ��#N���3su���P�`�R��:d�����؀\2��� ��P��2R���-�.
�������ɞ�C����e��������&������/^���)6X�v���i�q�-�zi��Q���&�UD�㚬yԌ!�1��Ͳ�ό��,A��𶞹��l��/D���̷�Ȝ{�U˅l�9�g&���Z�^ǿ"�\*2�\4(����Dj����/UU1che���	XD0����q�����X�lnI|���/�<����۱o�f��0gohܦ�S	;����<!e&�I���_�#8�px��J�j�6�&��0�[�`+N��	@�@^�H,6e�T�a&*$�@������E��s�X�Τ!��uΛ+6pr�/$9�N81 k�U�I���v��=��9	�{.�i�������~�%���x���g���mf/cE�;:C��x�"1`e���n��ln��ֆ���x�[MH�®T��S�`+���,A����?�8�H���Z۬��뒏UJ:� �w����6s|żB��v��D��ˣ�F�5^� ��p�����<#��ċu�X��[Nu��WQ��j���3���>9�+�&���$�:*�66��(�z�%蟚�t��9xZǂ�ke�l�{� ���$5*�~����aW���\��Y@�JY�J;L�5F ���$����c��m+�m'��r��G�ƴ����<�<���5��b`aY��[O�ۡ�ʛ�y�'z��PzP�8y���Ƿa�\�O��D#օs��qqoW6�����9���ǈk�t�y�f�;�������7�L��ց��`�FKE���ewU2,mV3S������5��D"j�v�!W`h^��V�]�l�1�Bj�8����Ɏ�i��t���E��'�ND���{���Qf1�>����V;�����7/���.� 0?	������~ ,n/v�6�/��{6����T�S�ha	�+m�}ac��Kf�86��m�2��|ނ�՞�&vd]�O��8���;YO-��?�?~]>[?4Ywp6� #���f',���=���4��99T�M���e��5��0����t�L8p"��Kp �������B逾�]o�7��*��ԺI�rx�(�V}����֥�����AɌ���t�S��xk� �e�H��>N�X�</��t1e��ShZ��;|Cp���	�DfI|O�*,���I�q8��U?
y��\.���|퇛N�հ��h���M������a��C�ԍ.���e	������FS���_�m��Wtѥ��k�H� rd��q�I�̈́�J,�~��f֝�e�+`r�7T �LʻM��#�b�Cs�#Lk�л��~7}2U��zZ'Lݬ��U¦K)t�jqi�h����]��G�j�L[Oð>���:RY1�Ф�*�좿j�=�7(%UHg� ��#��	�*�|��!s��uV�"��l�q�d	e��,-���
���Lc�	-p�
��1�2�Ӱ�Ѝ�g_�� �ձd��J��7)?ʃyDG�胊�8�JrS!��Jc��A|Xe���5̸g��;�D�����_����Ey4���ѻ$c����j'߮���G� �/������X��ɮ�R�G�b	��LL��._��%��~�`)�8��D�y ]F����$7�f ��$�?{��5�n�Z���;M�𯻲�|�P��b�܊m��8=@K��K`w�2��LTUPMW=�`���Œ�Jn��s?e�$��t�-��m\�	��C���͜˿L��=se��`!��;'\�FBg��y�jI������ɸ~��8��jiK���K�t�e_1�x�^��m�?Hc_��/��@�0�L��eIj�7InQ�����l `������p	�T)�ת�z櫠k��؛�	�bIfN��I����r��^�r����+g&cZT��x~08P!)�$ [X>R+�UQj7O�Uk�&OW�v�u[�;O�xI��R-�T(�_����i+��|m'`�67��B�0����9���odU�Iޕ�ݟ�	� ���g��mg�7�`G[�Q�r�r�!�(��������8�QͅE �x�_M�6H5�8�t�Ⱦ����]{q�mI�85�,���&	_�s�|{@ ��ԭGD�g�E؃u���ZR<?vD;��u�W�	}Jzܮ&ZH�>���s�	!�d+�O<E��V����_�Ie��v����9tK�L��T������of\�I"l����ދ����(o��zj`�q9i���	Ǖ���Sٮ3���'�
əw�$�4�jM�6��}��̨�ִ}v&֞jX�4��*8�0�0��dz�SXV��o�}��/o�ī���T��fT�2�@�;
���	�5l�g���K��e��l�Y����r7N�OPI���]{E����rnSwT���U��T��:��N��#�@��c��Ș��\S��$݋��.=x�u��+��d����F���D���#^���X6v�ׇ'�M����2K߫�X��I#��7�֊�sq����J�
��xr��D!��[��c�� Bpa�BiMX�p�k�uS��v,m�^�c�)]���C����Ά�ae�vp�S�i���)p����4��wtNΓ��s�&N1u�/v�$SI�Q�k��\#?T��u�B�#�җoTmΡkGv��o�[�R�m�(�`e��&��@Yc�`}`��9�U���v�E�Ee=/@'J��j��w3 �<���@~y|�Px��y�bg��B�8���Ȳmj�o��_�ҝ��w_#��ki|�*�P2���B�"�N��,N�y)dÚ��7ep�4Af����q.��.ڽ'?���(R�t��^.����q�'� �
�/�D��GJ��D����5����0=��{�l:C��xs_D�fG�������_\��R^���I�[Eõ�������r�����v���z����(���Q���tvղs"-CBg;��:ŒޙJ�����C[�p�$�v-�R�*Nhh�C �!��s�%ͤ���5J.�8dO����c:> 
(��}��r� �+(l����`W��$�-"W���y�(�X�����I(�3��o��z�y�8��U� g�����KJ"��؂w5dͨ��4�yM��04�AP�V�O�JP��D��W��9`�}9Gc�m� �X���ooEA0g��D�=��JA��`s����7��IŊ˯>E��!3H��eKB�7s,}���?�k�_�n��6��G�cS D��<~����!�KzJ1�4]X;l��"24�0��8�Se�Q?8���������ų+�e�k��tfW�Oe���9�@a�!�ޒpm:�D���Vjd�cs�$�3���-68��9ΌB:,��3/��T����aw��啧r�fה�0��/��K� ��쟊�8�,��T��"�C�a�ţyh!2�G�yi1\��z��N@i��Y�[�/OqH����go�/����ۉpl������y:$���C��B����1T��*���}w&�~܀@�IJ�7���E�d����iC���NR�8�i�q[��kg޴���Cu�Ǒ\�g@�{D���-�D6��bKtW�)e7��ۊ�������N�����~Q�9��Zd�yg�������7�py6�G�Q��/r-EL=3��k��N�mu�)�(�Zjs�Vc)ÖYQ����@��h���_�Y�G4UZQ�sX��1��¦(lZ��Q�j
�#?�q^��K	�Uh�o>�MT=.���..
��,=<�ɪcw,1����8��G3,R6�?
*� 9V�g���:!on�\���Q�S�y��݊U�d4s`WG��ڽX�J�|�ͣvA�4�X�@��������*�K���[��O�]�T��m��O��my�Z ����J����?�����c!l%k��E�)������>�k�*�ɪ��G���K�%�������+�\�:����Q!�r��3����q�bx�(a���}x,�^L�8̈́M��O���Vo���Μ��
<V�wq�/˥��୸��΄,��-�R�P*N���%l�:U�\pN_��mR�"�G�Z������_8GA$!�MR��v��W������fa^���lqx_�ʕ/���h��PXs�v�v3�CQtcz�N���"�⫏1K�"~"��p�������/�
ux�vDV��o֣��\J	GO�1�t��C[C�PN	,]~R�k�|4���>�w�����I�V�4�۽q#��^�a/� %�wW���KGʣ&�<��[�v�|ʺ�$O��sJf*E�gp�x�J�nD�6QhD���<LW9����f�}S�.�{ ��)f�ۘ��0��8kS`E�t��/OF�~�8S#A�%~��6�
"�3!�6Z�SS%:�}����� �'o5�XQ�"�Ơ�|�bȨ�h�y���� {#M�I��J9��"h�un6\��qP
��q�1=<y0����|�Q���fg�F�N�A�!ýq��.�/w�e�d=GY�I�8��h�hy���9e��A�)���P?�XG�Tf�0P�������{�ѓK�	Rm���`F�&�f��i�(�A_�$d%��$ۏ'�!�ب��l������.|����#rsAl��ǚO�����R�A��Ek�et��z�Q0��F7��0�EC@,�w���CӍ�/wa::&����s0�/��I[�:����s�L�YB�RI;��j+	^(v��t���H����!q��)�U2�G�����3<+��+�o?Y� *�o��5��.C�!�	��)�:�3�n���*S����v��[�vL�H��i�?�#�$����t�+�|�=t����}c�uN��⬢|�m��;~@;�c�	9y�:�59�TU��.�A�����룱��:�X�-2�����5���`�B
��==[Z��k<gO�eq�����L��^�$(l�8edEA?ĸ�1���	�sF��{�Z����|4Ƈ Z�T�>Ӽ�F�hE���%��G���|���Tȭ}Qw(�h���m�WX�?U� ��E��+Xͻ7Q+�^{=#�o�Pޛm���7a,ʒaw�?<�����6��=�Dz6�+��9-�*�+[�q�4D4�Jy�m�>��5�!�}��:ŕ���	�	��K>�	n��p#�j�5�h(8�3Ap��zK�������ɜ%�>۶	;Ղ�P��zj}����~�Ļ���)����V����P^<e���/���-�>	���q�M~�䱦*2�G��"̼S
�;��ç��h��i5|���8������S��Տ-#������F�ge�F-�����w��[b����Q� ��~�
P20���4�e�"w���%}�Z��	�g��N�GhG�Q�xo)\�`0
"7[	R *,�1�E�<��o���< �K��T����FO��Z�5�Ս*�.8ηˋ��E��A[��V>b�s��kk�)�H�qj] ��ik��~<�y�,�pX�d�=�%e�2?��jU�A�a��F �Z�I3� ��fj�����o��jQSwF�����R������@a��#�dI�����Jj���7��`Iq������Zs����5��1����~pg� ���~uR�>��������-������S�O�u�K���=4ϛ����ьI�>B<�>^�<�C����ì>����ܻH�|28�2ѣ�I;1K�j��L�cқz���Ɂf��u��.�n WBX4Z�v�_絰o_c�a:�hW���U��S���4~�W�B�����r�U"�KǁTa�:�/F�ee&*���
�Y�b�-�]�z U�M�������%ڣ]�\d܌6�Z�$�U���)��:��
���1.�ܓ?tD-�:�'{Ř=�޿�|}!>S���y8�lY���_VMP�]�w��l�Y�.J�H̐�#��#�ۨ���֞�lw�^U��αQ��f���Yu�e�@�ڧn��^�s,�����k��]n�H��9�~��*ΰr��`���8T�E"��Mշ^�~U\��R�	v�����}��\���jxx�Lw&�gVjW��y�]"����5�q7�`@<)�V?W0e�P1V��"�����4J���A��Q(К�BU�Z�(jH�q�rq#������@V�֎|ɥ�x��R��E����9�w$�g3+d(B�ʋ�-=�zыi��!$�s�s���94\4���?h8U�[!``�8�b�O\�鼥�p��,	�CJ}�n{L4�b�fC�䭼=f!y��+&=��*e�μwo���';6fV���M�׈�P��y�U>��~I�+��4�EN�ZEx4��R�f(��D�YtBDG52&!^r`�)�&�F��o�;�'�-�^K
~��:Y��<���sp0�F����,��g���)/�$#�f����0<�U������C��=4�.B�5~���ԄefY�Kp2d8P�|?@��EMM��r�׷3ㅔ5#�Q����=�z��Kú:τԡ	'�h�;�pB+,�W����#���-����k�i�(/�w�d���ȃ'Pk���o�AUmm��aR
2k�$�㷃%NV%ۓ�;(^M�Z�F��ƛV~Re.�ܘ��VD��ڭ��/���J�=�B'[�1��Z�7��������*eD��%�BLsM�b ��Љ�/����]tɗ�����zu%	Y\����G�~Ɲ3ct���#>�I����770���!
��ٷ#�+*@ș�H4����yW ��e|$	���~x��H�&*��X������	Ӌɉ�K:kr
��b���!�袼'x·�@^���e�>y�g~w�F���n�����
��M�VMK�l#�Kzm�*�̫w�;�Oj��{VZ�5V1��� @6�]_c��/p%7h1�SV��~,���_���:iťR&7(��������0��/I�N��a�?	W;����o+r��R�Ɓ3.�v7f�>1s��ڢ�̸M�-$�����:�;������e����m�����1=cR���
�ju�����)к�y������`��U��=�����5���y����k��{���_�g[]��scA�������5O���ӀM�D��y�$���:��dS 17���ti^�ˁG=�s~�b���[XP�U3����&�_̓iA��<ʸ�P�}anu @��O�AZ_�Fͮ���Uפ��Q�t����qIt���Nv�^�_x��P�֤DEe�"E��,
�a��L{��o>�fB���܅�l�� �$�V��~���^ܩ=$a{�Ͽ�w�A��6+�q1��ё���F�{�K�0��.�Y�L�f�ө37�.M�z�����t�0���m��1��`��a	���j�����/��dW�c;L�Wځ�ڎ� [S�������,[�C�NKͣ���v,[�x\F%�qw�i�ާn��.��2H&:2����kn*�1��?�KJ@.��/����Ğ]y���_aX:k��[EtX�8�a|`���F2[�/K36fW��h�8���C�tS��C2b��+:�`�l�Xfh�>�=�N(7AfXH�L#�6�U�/?�`G��D:�|�Nz2>u���^�̗�u�{p�/��gf_�
\6Rm ���F�J���}!�3����|쭅��=�^+�0&��Ͳp%6?��v�L����r�-#�� &��MsW�����Z�VUj��nG�N�r0P�|�U����Y�^�b"�T�������"V����(�b�!D��I�̴��C�d0X��\���P���X��1�A�x��Iu6��	�+v�l~�D�|�����ɳ�f�S�_�p���a�S?O��AIX�ӑ��؇����~�*�hv�E���>0�'�)�`�Ll���D�<tz�ßsr.��@�c*&���F��.��9~�mx��	l�LU�T�������!��h|6%2��ڞ�a�tOz�������%�DJ)��T{ݲq���0�O��KVi�u�Y>&%�����n�g��m ���6i��u�0R������_���p1�ZN�򪙞�\����"7�5�z��y���~m�i�6�Ɖj�X�_����#��L��]���J�6>�3c�S����q꒿��4�w�k
��f$��9n`�����2
ZǶ�B���}��M���Th/+k���,-���rQq)Mp��J_��Z��B��7���@l�I�S���B�;���F�5���j�	��C���x��M��5��׎/"����Dk#ԝe�XR-Ych�[jë?C�� !d�I��۫sy�/m�1���B�_='�[₨m�-H���R��>��ߠ�^���(��άn�[�²]紈�k�?�?g%u
�E>��WH�B�ck��s��X�eo���!��`����sJ���5�o�*�*�:*�a�U�X��p�-�y�F~M��D~�٢̓����<�����رR���K�pg~������x���?f�|љY%�"�tS��9O|���Z�X <�+��p���e���ud族M�����7�z4*�)�|Y�'nF����H���T�I��t��E���`�m�aߧ���q1&����'����T�o'�Er_M*)���@��"13�nrD�I����΁�ۺ�5fB� yw�0N1
 u���,�I̼ؽ�B?�92c9�K�S<� ��Ǹ|X�W�k��� �ͨ�h�� zS�3�/��3~�q��%G��R���چ-m0�kEg2X>@}NԖ�:� #y/��}O�CCΒ�G���t 	��a������o�`�<΁���֟��������~��o��{7��ib�H� A���ؑ�(�1�c_W�V|�ʐj�	�[nn
m��l8�-����-���dz�
���f= �z�>�����m�KQ`��+N��'��K\dҸ$#ivn�l�Fw�1�{��[�nPm�⣄IK�l���o\��N,N1F%a�ŵ~��a(�>{d�.ͪ?;����ONϬo*�T�lZ=�z x��y��ꥷ�I���P'�̮���8\>���o�5f�>+a�|�Dt<����x�,,pv� a(ĹՎ 7��*G��ZOE�O�'�%2�GW��-�	ie�u��8l*>6�{�Ϋ_��w)cR���MR��Y:a�!V��S����,0Q��Qwc�!ռ�4��p�*P��Xr���pw`��%��<�HB���HNW^�e��(;���DG+��|G����cKm�q��6ŗZ��]�p$,�|���5U���Lu�(�3���a����u.�� �;8te��h���$"�P��&T9.�`i4AӯAӳ�>(r�ڱ@B$��L\]�M����+��.�['+����N�a�uӹ؁*����[����1��U6�O�OXAS��h�X$k�ݮ�l��P1�|���
ݩq�FI�e>��l����v��n�{� ��.{C$6�y6FU�7k�y�z�V�s���;|�,8I^L�C>�������5P��T�_g�����+ޯ�t�KV�w�:���;H��ʥGQ*�{
�cu*IX��7±(����Zb�E���i?��]g^z0�?�ֲ��@v��p� 4��k��SZd�5�?wB�xb_��� 3���yn?kE��fM�)�>��F�����Ž�O��r�N�������
!h�S!�p33"Z"2�΂��r���[V�=��ǁ��)�0+m���┗x�%�ڂJL��9᪈�	$��
�)��QBY�'4Es���*��x5�%���k��>��9˦2C�=�@�I;Uªj8	������(�J����:{^QW�v�o��49�|Ր-�u�4	!ХtkDN�#����¥-1���`�HD��ML���~���)�'gy�uc�m�k����섄7�B.����m�����[/��=��YiUڛ
��f�ܛ#�Jz������y��V=A��@�D�&���Y�3�e�'��� Tb�woNTc����g��7�=p�q�&�r�ԇLFPl�hKr�e+Ҙd�5�\s݁U�H���Y��[����ϐ��UՆ�"x�|�vٔ��B<|ye��,/=.���X�F�;�7f��l�����@ޕ����0�/^d�Z��'�j����&�|>�6��>�[;�C�Q����sMZ��kr��<���DBr��(7�d�>��xտ�t�M�g;͸�lO*F�k�k�_�e�4��1��I{�`;�6�$Uv f<q:o�k�|�/1S�O���Z'{��i���n�����ހaL�_e�`�d�"c����܂����l,x8;O����h!/�|B�W}��ȵEұF~f&��]ڴ,��\�ܦRV���uD�{����5��yz��}f�#z��R�̷��N���c)�}�|�+A�q�dm��wP�'�>�3�LK����F9��F������$�o�J�̝�E/�_5�|?���Q0Y`E�z�f�UL��9�f���ʿ8��W�����l2�s�>]�x�Ad���8|眑�������r���K�:��( ��f�ܽ����>@J'���
��Zf-�`�̠y��J���Oz��u���<��\�F��@�/<�ǖ�-�a�ht��ݩ�ڢ^.��:y�;G��HS�6bc��⤋=�J�����i�Y|��wR a=�+;zAR�a���E���t_�G�M���doj��̯Lir�c ������Ω��7ڭ�*���U�ϝ�E
Ԉ���i��Nl�6�Y�:4�[�\b'�m���Ӥ ���"2�ɋE6���=a�'cb�?�鋍�]�_�����X� ��m���5���ɺ���;O��5�6��~�Ԇ�Wĩ]���f�2�H�$?�=�/��$�`���z{�+E(e��aLͣS<�D�qCWT�ʈ�
[k�wu_~�Q��
v�O�vE}��E.���txR��Ԝ��	�=��X�[n&��.8>���$���㸊�!� 峹̥i�a}7��'a�-c�va��P�
��u�aY�җ�,~û$�?L�y�~��Nf W��U�ځk�/���I���V6%�1Ҿ�Keŕwo ��˭��������d�P�h7r��?��{yJ`k�e��aLW*1՜(��,3EW8��2ܝZ���D���D+i�C��D��86˹��
tS�.�kΎ	�O�%TT~նA�=d�i��FV�#(C��WJ�!�l���Oޖ��cCr�S9����傋���E{]D-�Q�㖚��
`���Q�:�U �۾��݀o �13΀ic.����x�����@�>��&�ƪ�d`��;J<$�?ͦG�w���e(P��|�1N���O�;�'�#�]j(h���H���p$'�]e	M�T���
���|����/�Up,\�qL���|�-3��QUNQ�J�*v�j{z�L�;-h�
�fC�� Fp����z��5�U�&�͟h�Yyg�E3B�X� +������.��ͳ�,m��DӍ��c_<��i�:����(/�@2��<�ش(���^�+|5��J�Ԉn�1�@����*C`�Q|@���/��zN�uD�k�Or	"�/{ߤ"g�$%DK�R���ݡ�i�c!Մq"/oi���%�w&\U��:��-a�� "���(�g������8�W�خ�b���r�龃��WA�}V��qu�'t������O���%��g/�),�����9���|l��R%���Lă^����cKOx�J��l�J�I�z�-�7y�{��S�#HVϡ�	�}k$	3a����JiI+.V�y�2[ �'v��+��aڦ���~��&� <M��<�H�����4���TW(E�#x>9 �H�`�@�\�pV�'�8�H�ɵ����d�(���%$��t+��*ՏO�T��V���b�wih�/:I����`G8(D'v(����JKi�+�s�D�k��\ �v����*�����)Қ�@v�!�3�~�,g%�6�WRƿ�臀��-zd{�j��N�;��OW�����ltbd�2H�J���'�~d����<�
��6޻
�.�li!�|Ѣa��
߇��C�?�R�iP��Zy�],7Ѡ��H�تI�E{�)��,p�-541 6K�mR��b�����!�55UxD�cgZ�M�O�\�;mL$*�����[�=a��w�j�SҐ�M�bN�6�O6��F�B�3�������_D�
���C�xd�'��>�ν��A�������߈�+0�N@�Ъaο�acEug�Z ԽX�Ml!]U�l������1�Il�#��B�t������~��~ ���V�t=qs��_�Z���-S9k�YJ��gΛlB>G�^�ѴawT���sI��/猆4ȥ��D|�a�Y7=��}>}����[�w����Qͽ�R�ڗ�3�Z]��F�]-���D&vE\%�S�QP���Q��K�ʅ��+c,L.[� �,x�1-f9���.�'c!{l��΀��):v�.p�L�	|97_u>�����Y���H�V��hXM� ��L��JU�K�M�jI�+;� �.M�����o��]����tI�M��-!��h
�b�n��
~����T�'
��빂��*4^�\�����M)NZ����K�}�������o[a��
 ��ŗs߹N,G��uW���A�-�i�v� ������Y�����IV~y
�]�i^��m����?�e�ڣ������5W�KF�Ӱ��f��
K}��;��H�x�6q%y�.Ta[eΫQ5Î(W�zc��L���~�0�A����g?�<��*跤�����v���D�ܖ]���y��z������>���D"[X�>y��`1I�Ly��y}�=˻�����Oj+�`L�z�)[�>~u�m�r�<�N�����;�^�f�N�=s��?כY7��r�Z-x�@�����(��]��5��7�JVF�j/�8�ސ�cO�z����5����h҄B�j>7�B
}�	��z ��l�6Y��:< ��n��ث�y���ب�A<M`|�/�W��7rE���hϹ��?�QN���t@@#Ϸx�h�`7��kt��c2�]�h:��L���^Ga��]��{9��vTW�{e����t��{�ӳ�k\5'%- ���>Tw����C̊ȝ�J|A�L�ϗ���P�rV�}Ǩ�|���0/T�t�-ņm-��q�S`��`��sZ c�}��6}����iI��%ޔ�"�G*��ˢv80ep�sN� �M�uU�g8�E�|7���H<|y��K�O�.�VO#O���p�Z�v��f���c��9tJ�(f@��w��C��9���z�{i
#��2(M3)�R���8���BM�ر�,ɳ*.5��ޞ�oܐ1�S��?����:J0AY��Ķ�Q�i�u�y|`#�b ��I�pq��n��M�)��TMUj8 B���7�x*�_�J�^���rY�PfV>���ɵ�N��'�ŀ���B�m�o�·���N��Mÿ�Ԗ\ $�`}"��|�h���2���9~f��
�%��0���Ȑ�q8����$5\�c�����Jzi�6v�w�h��i��z�_,��o��3k�/�w��Wv��l�����t[�������:��z��=�\*a�`|�Vf��6�;�B�h�b@�^9F��?�7���`KJ�%�w/�u?ӝu/�z�}�'�AO�nGA{��`x�F�F�_�ػ,������'Up�2b�-�� yr5��ԴJ�!a�)��	��n���S���D�`j��˞�I?���1�]�pL���9_���p:�-*��������TV�O���Vy�s��r;o\��������>�B����Cx���Ⅽ|�w�t��F��si%��מּ�ƺ��"}"b	����eqi�����bxQ�g�<�����h\0�f)��J{	�XsϷ�&�r=��ά#	K�c1y���e�*�:�P���kv��T�)�$>bR���Ս��\�§�RS+����|�s�����WWh_;:���M'QR���7]�5.|�05KII�t��鐶:��l D�@��i#(��_-��mUBV�����ɾ�g��B��'��Һ�9:�`��9�9�<��k�����x�~�5
�$���xvP\�RJz���'�0P�
 <�͈�S�G��k�jh�q)Y����Ӌ5�Ep�W�M���P~&��D!)�R�rF�Dսʲ]c���bN}��V�8ð5�:�j�ܿ���^��J�YǨ�*!#�4�>�
�%��!�fd� A�=B�0!u���r��Kk������_���@��� '���P��';
�᳙ˈ���h�ϫ�@0%���2�FX�R^FW��E���t�$���1������L��f�==���o�>��ި,��3=:gV���x*=��A^ m4����{ p���]&t�x&��i�ג���:������	���k��l��V\,Q���Ð��J�PYנ���<�B�m�I�2�U�u��2�8%'�7����)�$��Qi�W�����Z�hE������)v[`�UL��wmr|��>5�$�� ���e����
͕`��	UAr�i������2���.���9���J;+<<Gs�o䇒��+oܼQ�����$?��򖟮WP�z<)Y�g����=�Z�yL;��9�_˻&κ� Rm�������V�4�����Y>���k��`�w��0�>
U���SxRc�	?��W���S4t�)f�x�h�f7�s}H���
S�F�R!��1�u���3ִk�{30 [��1~�J�-���5�M�<�>e��Ď���_
��u��P�l���u9��L����Ǉ�D����6{`TO��\g��,QV�P3Cm]��s�	�=`p���/�o���LΗ�O���sp��h�W�����3�vsiA9�y�17�*����Y�=l��c�L^7���	oŃr8��?$��R���Bb~�r*�fֈ�hQ{zN4YV!~�R(��q9WyeH����ٍ��Εw�;�6o��$y��eka00MH<n�X�+��)�:m�G7��ϐ����Z�J��,����m�����<VV�u�}N�������P�]�gon��<p;�켂�ַ�zv�b�_�kY,��^8ڀcwf���c4�^'��Rq^���>ȫ��_�s���;��>@D$��v�a�U;$e��3�J�{��.���s:K�}эv
B�t@yi������h������������Ki�EPh,�O��x��;�<����,rC;�;O NP��=*=�Fh��s�K�ӓ�B��	]�Y �<�<�]��_;�_y�[�1麫���`��u�sn�dG��Rfl1�-��\�H�y�CA��\n�����e�����'�*q���#�a�I�=+N��-��h\��8�#ьdc�۶>�	�<�IT`Bf�f���8Q�Q]!��]�ɫ�Y�0���&IO�?����In�d�LW���ȷ�����kX�B�C�\@݂��S��ʓˁ�6v��袛���f�)�7j�c���P��˃�"2��2ji�7Z�G�T����T��7��b~R����j��4�;�����g�o�������e<�ua|�A%ȜCg���;��5i龰��ړ�bֽX(?lmY{<\�	z���{�ɽ�P��tֆ}e�*+�.��Y>)NuC�}w����� ��6Oo^+�y�>���Q���^�
�g<�n��AW�����ܹ���C��Czp���=���I�2f�ФDz���sn�[+
�h`��5�ED
sc�bk0F�	���Ƚ�@~V4~{��.��(Y��>�مk/[.�H�'�2sS�p�HaW%iYp���y�E9��"�8�� ���7��~�M:	&cgK�T8���t3m�Ej�|��@�:t����zgKWj�T�klދ�v��ͫ�:U��=9{ْ�?<�D��W�Z�K9��A=�Ϋ��Y�Tn�P���5�k�1s��j��<���l7+>�����P7��X0zy�_6�+k������3���/�H^P�/��.T��>X�b ���?lٱ�ܒ���(���(GUvod�0�(���B�2����!�S�l�[r�����T��Ң��HRX�k��D`�%Z�Fȷm5�f�!=�W�ƪ��92�Ru�IE�H\V���t���-���9<�A�M4�J`��h�EC�l�:m$��*qW�"�QR��`�1dO�=�5�~q�w�a��IE�y�u-n�:���̣�����k�ަ�p^z�⚟��x�t�6eg���N,c�ha
���ַ��]�)֓L�>�jv c`��}ơal��
�HX�������N'H�g����XT�Pj���?_%?�k�:�:�
�
�1���� bv.���J�ܔ׈	r"���?SA�h�>!)�8���f'e�u��c|�3����
Ȃ�z�j��BAeT�F�"�EՈ5��;?��S���L���.�
q~
���"ɮ8��JU��V|$
��)��s��8��g �7����!�޲b�L#�%��������y�O]�� Z(��a���j5f1V�[��i��E:r /4�l,_��>8��n#���AP������>��D���'�,y���Kɻ�����pn�	�dZ���,�I�%?�p/~k��p9��=���ثk��y��1>�xeB�ꀧ�c0H����3��R���n|�Z�
K����b�4O�S����"��/`d�*��>F��E<�iZ��s�{$ˆ��D�r��T�����Fg��`炾Qg��-0}owC�"u�kt&b8U�S=du	 �~�j]�",}}Ң]81�� ���l?���t����
�Us(�X32�ӈ)�-NKOV��9]����`14'ۻ���,k},��d����6�C�K�FbJgD����q=�6sǹ)���t[�f�*�(-f���k�x�^7�鿞p���g��N��%bЅ�m8���&�!�n�#I�mr�V�(E�TbA����S�/q�$�&��.�Q�p�^��zw���19���S9�1���B��쇺&@H�p�Yf���"҆bJ�!�¹y�=W]�>�"h+�H��m�(�cHwv��hF)Jp;�)��؍q��S���Xg��o삛]GU�|��Ftt-��o򀥼���AϞ$�!	��*}�'�%6Wht?�f��<�4��.�U+��޷���fۗ��+��B\���IL�'X�%��ǲ˄ 8 %e����0]5� � �)6SP(*�D/����c�F�x}R�PNKط���"RS�i.���}�ōs���$�4'�B֓�J_!�:a۳;&-���("���J���t-S�����Ι(Bw�Єyâ]F�͈���]��u�Gu�VykB	��,�į�x:�4��g�9��x�<Xbz��;C@u6�E��ˉ���e��I��V\���)�{�&����{�ue�ů��k�r䫕l�f��w^��@X݇����B�`h�Dg�:|��,0����Y`�{F�V@�/(}���f�F[�F���>;btb�@��qraS��W��>��Sq�\�5��X$���/�w�Ճ��ral��3X���֢����Q��$YY�.�b<ݦ>�H)��d-y�@��ƒ�ë/�a$�8e��^�D3�R�4벤>[���a3̒@n3!¡#4��5m�J�.$%z��"�����*{��t��N��� d'W�mq�
�ۘ���N�yc�岘���Q�E�%��`cWy��UꛑR��D��+�:��jL�Ӯ���ٰ���/�5���Hy�m�?�7�c�:k�紬+�tR7��1�����,W���WI�Y��p������$��cb�ư��0�l&�t��(es��z�1��;y°�p��u��V#���_�y�`a@e�J�Y0|�|R���Uzz�d�'��H�i���z��=���}KE�.���0�� ��å3�?��`�<$]3�3��ɸ����z��Kk�5���aK��B���y�G�[�/?�	ܤ�^ ��=%^p�~%��k�o�l% ���hc��ጋq�� ��^V�/�[�%ͱ�Ū9��� 闧�l�%-i����?��d��F�^l�Z��!&�ۘ��h>�G��]x���8�r�GWo����L�uԃ��g�u�տe��CD9�3I?J�j��q1���s��w�Ҡ�qh6.�8�#�V����fq��[��>)GDU'h_�[4/+�Ɍ�ܡ&\��9{��/��H�Dv��+�x�d�������~h��W���۔}�ZO8|��w���`v�{돆�^��XA��9T���l!޸ �����k �������K=x�T�����L�&b-Av��ia��X���ݤ�x>��K�������*%�'"�S��.�tf�����s��X�-�� ����c�vD��g���~�$����� ��!W����r�1+ɼM��!���~|���?���	TC�,���|���GcW�pe�תf��nS�D��B ��T���tX���#���l�d��k�_�#��ѩ蝭�X���,�4�L��'��	F��e.��;�I _��(N�I���`
����'��ʵS��=��?�-o9b�,?J豷���m�h�o��߱l�o��-�6���?�tV�<�>q����JdXO>H k�%��{.�&�X��}�%�E{q:i<��O�lZ� PDHv���y�r�_��0�(2�� e��,��F"�8�ȍ��[�Rjx#�m�#����W��qNnR�g�l^�⃉Q�͓C�=����P*ᖀdI<n(��g� �5��[eq)�b����?iM'�V�7{�ɝ-ŧ���� rd:�d�JH�6f!����4�Y���~=��(�@����؉�PL�Golf���wf魳Ƚn8%��'���^g,E`����1uʚ�Wk�����Ѝ����r�� F��1ŒH���qgP-A<��F�0�]��Y�D��L���{���hF:uC@��X-[hz�O�.����{윣|�	w<F�����b��qʭ�m�7���q�� R�S51�H%[��>�?nx�o9JUP�'��u-L�HV��*��(JVI ��R�m�0�\�C#2�!;��O|4�։�cc�������/�=���g3ϊNxMMf�iTI ��2\��-) D���4r�e@w=\��b�xs��܇o\�t�(������WW��J��iΟ������|��O����`�1	<53����/E�b�)���U��cL��R���L�Ǚ:���݅);l(�r+�s,j^QQ�������0,��$���%nж�:���x�B��n1���5){��Z�S8g��74�M�{aL�#�No��p�!$!O�J��OL;�
:2���^��� h����H�Io�(vt��e
��z1�&��!G�s	D.�x/K#!i�B��WCbm.E"���7F:���k[{�����j@J̏O��5��Ǿ�IŚ�WF�Ym�&`ۅuo�m�:��;�QPJD�*\��L����!��$�)D �2���q�rU�l���Vh� �Ȃ��ӝ�1��2���F�Ő��)_U�2��+��M��~e1���)��x�c�X�;rS�i�!`���،����]�p�2m}�^����a�Ļ�_���3&IW��`P�ZW���oE�>�����\�Қ(̕y�09�Kê��˘ޤ^��Rgڂ�����Y�\�D��8���&c�3iYrtf��@Al�t��op�ꀀ�k>a��ʌ�,ьP��:
׉��Y�}�lF�O7(	�'l����]Q*~R���D��=���u��3�A���x�?'�W
@�Hk��M���7؄U�+�q_��D�a�"G�� Ԥ��Y�"<��O���q5^��q}�,U*�0����9�҆|Ի�H�fZ
ŉ.�,2d�#�Xί0�^g������钲�
�)5Wx5E�|Q�YÅ*u�
 2�sz��!��6��i�	�v�&<$��U� [���e7�����E8�	�-.:�O}Cfm���8�y�t�S8~I=|���{�uYXq�걑�@f2�7�u��a;��K�ה��}Q�M�*º[<�f�<�V�����ߙx�j4�"�b�#(���=��1]%^�:j��?�,Qţ�'h����T�J0 ԡ����ϯ�ְ��? ��^��uj_*N2HaVG�Ƶ�A�ȯ\�W=!555dq��)�ۻF�-�hT$�b=1�* ��߇`��㨶mI�]�ٞ8].�o��!�o�b��-ߪ���Ւ�A�54|5����19^�b�B3D���Qx����J.�+�BR��M �X{�Dj����
w�J�c55��{�Q~�Aͺ��~���f�g�Z�C���[-CNC�5�=�� AkyK"�a�ͩ\l�-()_)�c�Wg8$�~�Iω�!��u��׊�-��X,6��U��|�� �E�*�S�˰�lt�`�8�=�	���ʽ ��z���B�bI�I��fx��gWZGOrD�ς�8YW͎R ��C{&M]�i��>Go��t�j�|����L�Ts�^1��}�\�i��L�˵h@�=�9��»�f��_����}����p���E�H�|���;�FE4ra[Yl�U���}&�kB��~�uA٦񳹡�8ke�� v&�gߤ\K��R�x����;Ř�-��)�ő��At��M)�R��>
��.��Ņ]}�L ��P������{l^�b].o���ō:[LLh�
��D)'�����RE7:Wgf�|X4��K��Yཱྀ�w>j�4�եc����[�i��	u|Mj8��o����ky�F(�-��m�3�%�e ��3�+�a��ރhb�8iK�)ߖA��	Z�{s�ʊa�#���7S'2�`?8EC������ۊDI�kqn���C,짾R�$���Ѥ=����z?��̦�����U�N���;ӝ�{!�lE�t����]�����	��2&�������F^�im��V��c�=W��J7� �x
#���%i�|�O�~#�XE��� �����\�R,��k@��
K%�M+�HǢqm�ѹ�m�� ���C�0摭u�-e��  B�\�߲is���҅�_�'ʟ�q
�9[�'�FL�F9��q�\D�vNOl���?��O�z�� lj�T�J�jm�����nm����_D���ˣY��nS�+��"��z ʁ<�Cu�h�A�=�jz�z�z;6�h�h����(0$t)>Z��
�E�?)ș�������}�c��I�,�/��'��gkr�6��_ɩ��� 8!b�*aQ[���S8<�g"S(�w�W�$�ց���],*���u��F|��B�c�����#���>z��� �]��l���mg���tf?E9��d�0��e]<�=YRKf`�����/ϙ�8M���;����zA��F;kY�a��U�-���(Of&�ɠn�6�����v�j�� �*]��#�m���n.ōG��ƎJ6!y@D2���^J��bq��;G�d��m�h�T �n��e��PRٟS�v�NQ�yɭ�rO/��*r�^��Z�}?�䠋��h�':*G���!΍/n��J(��m��ؐo�����{Ww��γ3�P\����]��W9fO.FV�qB�_��?��@vmd���o�Kӱ]���\F�J!������v�8���H���o�pNL�u��)��x�w��n1Qx������E�>J�zG4�2Vx��.X��
��9�|�;9-�Os�y�ۚ�l��զ�|�LH�Ⱥ��I���s��"��{����q�����S���������-�����WE{�
�KN�}5���Y@'��s�RW�Ц�b�W#��-�O�r6�w�Z*�{W�0�y-72��X�Y�bJk1
��Z7�&ٌobM������j��u�尤�IKП�����dKL���tO��G�^��*��ah��g��mo��7���I�����u�RWGƶ����rZ�_7��ޫ���:	���1��t I'�Cc���[�`%�r����N���vEa�ә:o%��4>���]�.Z���f)�m�˿��6J1��h�;��p��Q��GP<������uCLk��K<�m��V;P�_���$����)#��W���X�5W�`�P�h��/Ja���͚�����2�	GW2���ucd�$b�%��WO���:���1�c֪W	���o����p8GJ�/3NG��<�>gTV�=��$��k^��i7��ZӋ�ac|��v�CY��9�m�\��O7 �	���M���z��e���x���at:
�b��*�C�F���C�U�c�0�4СX��H�?|�RA�X	�c�˳��
�i)	��|T�����t@`!��xI�/��]�X0#{!�P<|I��P��KI6Z����j�m&�f;(�|�n.��e��:��	�k�A3���߽���3�����
������j[�=Ks���6E�ý}��_ҍ���Ԭ!�sJ�,yg���(9e�u��:}Ċ�ع�3�J�Qb�40G��Ɣ�9um�H+(�یt�?�6湳UAY$�V���ƿ�͸�kuᠬo����*e��Н&9Ш�M�c�I{	=&���z��:t��H��%~��-
�N��z'�Ì�Hü�[[ǥ`ݘQA�5�Թ�j�:0�3|lfxI�Ji{Vv@YH��=_*�J��qd׫6]3cߓra]����$�
Az��͞��7u�%DOR�Ԉ�J��9�h�^2�V:(U��`�����(_�6v*P�11n�}�x��w#Z����5tn#�R�X��3�����%�M�3�iMxFS�qb�8W�D�������|y��s ks96��|�k��'N2�O�`7�Z0�7�ޡ��!�I��}Ϯ J7�(�?�H��6fe��GOZ��@@�����7�Z�� ��X@��%>��Ssd���7J�j��Y��y��`�����C�^<W{�W�6�G��r��@"�:��;�M�p������'����L��
E')u>&8�ڍX�힯]@�<Ғd�Q����q܋�L�����y��|V>B#,~�7M柢|lr�*Sg;�>��*�"�������ھD�7�e�2R��;��y�w�5�l�z�n�&m&m�i�v����)�v����PN��`���#��E7�<=�Q���К5��]g�lx��8HI�_L��C�Zt�r��3���d$���o��S= ���*��S3ݹ� ��Wg᦭2�O����&�� ������2h�x���g]�cG�/�E��GE�	>�8�H�/��T�,x;c�z�1�-#�#4*J���O[}R�����	sF"��J8H!�׃�'�^�	�ڜ���xc�[��7	}�P�I�o������I���Ó�H/� �/L�b���a2�=Q���^VP��B,$p����/s�ݠ�
d!tM�� �f5	�M���w���#>A���HC��A�͎�M��-����\���n#�N������׹Xi4���d�l�]�,L=�/P�޲�Hw/�m��	��ĩ�'�����؂vA�����ܨA�n+*p��bcMu�.M�}�M��ί��`���G��P�k�-���$��J08Џ瘌���fN���%v�  ��!Juu@l�}A�o�-f�#>y�0���1Ot��&�&�Or�z��DE��jYAF*-�� A��aV��T�C�'��J}�ys7PSX�M��9���X��@��M����������AڗX%�8n���{@RB����Yh�a�y�d" ��G�5�f9܍�HX�r�Waqؒe�f �$B����ܙz��g1������E����[�G8Ib0,����(>f�|h�D5�����8��b��j}O�s��@�?�4Rur�ej�da�j�S���mX�]D5�2�K��!C���d�����s ,������D�Ң�2}�=ۺU��}���>`4A(\Ϋ����3ˇ�΀/]�G�������6^K��n0��s	���*x�&�)�C֚��Y"H�E!����Y5��렩y̯4�����<�x����k�M07!��
�{���R֐��!��ۿ��; ]͏	v 4cz<��.�Dk��]D�����R=��蔞C[���|�D���ʭ�3�
l/V��>�ԁ�Bp�9�0�p�����ը|����5�G��W�JX~�)w�U�F��N���X�^������Ձ�7����f�ݴ0��lh}��)=�T�c��.����1�o)�^�3b�v%���ae�콒]1pu<��o�;gЪ��N`�G�_n��q@��Z R��>#��ay�{Z� �Y�w�����VlY�I�k�e��;����Á��	4RG�j;�z�x�9��PMo��{�[v�0�Wۯa	jِ��(Z(�	�:x"�al�3ۆp�h�"b�n��@+��r�*��ǅ�X�+�#�{Ǻ��GU�|A$U�g{�*�/�Ҋ�ٺT_���l���N��c�p��ن�-���#�1]��Ѷ4�4�����07�����-��'Ki��&���1W�Eky�E߅r��S��\Dl`�U�]_�wu+�#�En3�.�
����h+��>~���[��*�	~4��1�-�n�����J. �i1��mT>�M����B��ƛ9��P���*������-���s�^y;;��Ubَ<��m����?��+K�+{�gCqae�>�?-�_�>��.����^j)�5z�#"ф�=���ó��H�{�[u���d"5Rnb�������K��=Uy���8��U�5Q���#�@d�2s:�]2�]�o^֞1�6~Ġ"%e�WA��z�F�v�+[Y%��%��@��Xdb�|�8BRg�aʞGU�L��W-��Z97�KQ#�H���"���Ƶ0&#��Tv�GI��gU{$����WgT�H���sd������cn!�����tB���$}�E����2T�@����Fq�T6��B������(UY(���w8�'���(��T�K�nO�-7܍3Ў7��yN��ڰ�t�<Y٫D���T���)n����y���(1OlX�ȫګ#v�v�8$��ECĵJ��p�( d����
:��U��v���Y������P SV�w-:�<?�{���L��B�e!�%�Jq'�x-k������"���j3�KW"�goϷQJ]�@�.|tj��\.$b��.%��.��P���$	�R�R��~�D��*[�),a�\vz�mW�w����@uۻ5�M$
wʛ�wy�;��c��k�6!��t�	i�3��pXnT?����y��%y��M�Bm��*Ƞ]ʩ�v��,����v��l1�d+��m�(���b��?��R���Ƀ_!'�i��5���d�H
%�� %"�6"�%ME��g�ɼ���R�]����W;��y��M����y��b�,5���s�������oyUzu���TU���O��%o��eq;��^�������G�\�I�Ep�"�_��8x�&��b�R�;�]6�D�z�@��-���l��lG}Z(y�;$	}��{����%��A*X/�&$d�I��WO��,}�KD@��ъ>	��U꧂���;���5d�V��������%i��*ú��Ii��s�}�0v ���C���I�)��JZ�N�Q�k�KݞW�
� �U=)��F�n��j%4��+$H�:��=q5�j8��W ��A��X}�
9k� �R�%|��2�#���:z4�m϶ˮ�8�q��:s[QSU�	y�uQ���+����H�z��ү���y3R%���H���r���\y�� �YLG���cQ_���� E �d����t��Y=��'�u�b����*�]��g7?��_4���!^�W}8>��-��v��F�
��MP��ǣ\C��&���0Ā�`ޣL�m'.�հ��k�81d�,�
5�JG\/tSۢ����<��a�+��e��
}�0aA{��"�ӼJ��W�e�x(�m;,���ҐΎ0����k���l?w+����q���6��y��)����O����7 ���F'�fׇ*���L����+q�so�E�bԌ��(�eL��I��%�~��;=T�7�E��vģf��Qob���1����>���w��	�;|��@$e�@Pz�pVH��4u5����H,���.oM������3�"�(�9M�����M�6��u+e:����-�Qw�����J�)}u�'�A��ؚ8 Dd�f�]���u�7�/u���vQ��P@���I�AD���:N�'������ 	�#/C�� !�i��{^�ERdB���F{&6����MD�7�,�a��ix"b�[H�i-�3�S�d-�K�Mڿ.���7El�o[��#�|-ЕE�w/�@�>�Iҗ�i���[���k}o>��6�q��'A��T64�cG���d\���Ih�@w� ad8`F�t��g ���Q��k�Xdq�����e����Y2%n�U:�K'NZ�����j9r�9�y�=tEқ�"�GขS�F����ԊC���?�9�xi�Pw�L�:��e:-n+�i���=W)�h��<c�͟9� ��&�w<�zƦӑ��b8�������Z�o=[[��4�*���#3��S�,_ Q��{��V"<����0��؉�Il���Y����E-$.��S�Z�"��c�~q��A%��5�X[	���\>�OF�E0g����2(��$t� BF	�&�μ�3P��P�B̆������U�r�&�m�w�������-�Կ��2ܬ}#-Fz	���A�e��R��&}������,��}�]��Q�a�1����V�qm�,1S���RL"�C
S�}�����Ul���k�����Ɣsz���A��X��!����Y�����-�Vt�d3%N1T'2���FM�Ӿ3�-"�@9-?Ql[`���^q�� b��"�X���Ϗ�#��߻��Ol3|�Ĳ_�=Wӄ��E��Q��ux|m:�m�BɅx!���kI�9�h]f	�w���.� ���6s��%ـ�r��h��,��7��Ij��`��55G��-,���P��h��ƫ\�>�����cZ	��,��m[�7����a���&�H[@��rL�&S�3���ȹoūd��E�Ә,�j4/X~��'{C����b�� ����=�����r�S��S˕�i@@�T?Tw Z����IK/!w�D���c��O���4�Q�`\�^b�;P���C�Z�j��˪�,ӌl_�L�-:�c��w݃3����D������Sy=�=��G�AhB�%'�4�-WT��6�vο+��(vȈ��02�����69�=�1
HIHQ�X��2[P&���@��Lk9��_q?�4 b[��=��O���˿Մ���Y���qlE�˳���$�KJO����K6���XT�b���2�c�Ӏ��[�L�{��ô6�h��A���F(2f�g��1̜�;�����!��B
£PY�T��^c�m�H�������!��m����_��p�E#��7i���͗/C,��4X �w�Mr�j��I�_���RF����N� �W _9.\���5��O���I��9ߩ! �f�	���<�fs��]�8���K�����[ޓҏ�R�2�H��A�:xy��-�ssi;�[�2s��67����H]�:�@�"����iE�M�[֞��&��Ƞ~�ql���;�X�-��w��k��b��.�
9v����5�Eh�P�6T"RD��e���=�Q�)juֲ	ܛV�� T������G��Hb	HS��.�z�X�F;�ߒ{c3�H�C~�7��R�Ѭ�]���"���j��������"X�11�^G�w�Vu��Z�9+���{ ��x}P-�X�j�Y6�����F���}\��G�_�~����M�H�LcI��׌ˬ��k�i�4��A[���+3�5j��D��3�����Z�FGI��d�{R�6M�O$�s���U^%��JH�z0I;��J�=z�dF���&��K��>�NtB��V├w��}�d��1�˼��,��о/�P v�M���h@?���ó��5�������r�%�G�Q��.�٦���ޓeT��B��!��S�6���X����a� �H�Nڅ�,_'4����hV1�n�s�)K|����7n�@-q�!22���"4L^T�s4�-�K� �Z�bE�xG�,��E�U>����J�)������*A�Z��aF;h���J�{'eʉD��>w�@�%����˓?Q��RQ��?K y�s�ɓ:oWاC���"��R�=�Ι���j}�`������:�}r^�R)�~&s��z�I�m��E�F�oi��r��B0�2�ˠ$��b�*R\Z��[�	�sBqC�<bf�nA
�"�^wQ�l)�J��\~U�mȠ����u��Q��t���wx��?s,��+�-�Adw#ZN{�Xޣ9�R��X׆���w]�J��ɰ[!��hЈ־�FH��m�7'�b���<������k��0�����0�������=�D��T��~ރ��m;$ګ�sh��4榦\d�O��Gx�fHBoGSl4���;}�s
g٦���R�b��D.��_l���:�}��xjB'0)���	���2f��hj�FџO�N���r�7��y�Y�.�f��z��*P�@i���
M��e���/Oo��r�L!�y\�i>�����H���#�#�<�CQǀ��'z�sr�(z�'J�GuBw�q+��;Í�Km�Nb�I���q[�w��j����E�fޚsGjܧ��o�Yg�"CV�U{e5��z?8�Z�Ҥ'��c7U�5��9���HAh�hI��{�`[,
��[�p�/N�L5P��^�S��}0�L/(-�.�7�MKKF����y���n�Ʀ��:1.� Ba���������;^��,�����ᨈ
�:��+�}?�d���7d�Z�;����64�����Ga�6����A|�*͊�zs2R���>e��v��^�a4s��r���Q�dQ(욐~ܖ���]L\�
�OK�/�U���o<�b#-+K�U�;��Ƙ�"X�����,�=��$%m@�6Wj7g;h�	���� k�6q�e��QZ���W]!kjy�+�O���ή��DMU�-q�|DQc0���`��
�V�c��5�!���q�����4zv��i���T���ڳ�DW�@zb�����d�� =�R���
���Or�uB pڞT�˸���9��h�N��\r&�t#^���}�bƜPG�� Ϊ�W��ECg{_��&i֡�*f��V�^U��{��?2NQ��=�-�l��m�9�m"{�_"a�7^Ȅʩ�-�c6<�[����Xu�� 	g�eG}ughZQY�?����y%���n�1:�T�a1v��_j�Ѭw,��Ȯ�����ͫ{a��޸W��':j���}�k�,��ӏ��խ��h�?���{4���,1'E��!_�U؀�op�Q�`"u�P�NM�|FS��	Y�\R[�
�t/�뻨VoΕ
;�}�"d.�簔3v�W�r���k ��I�{�貗��[sD`�KO��_�w�#�����f��IP�\�
���O�դf'u�b)sݍ���}ɶ(n3_�W�oq̕�%gܧ���&���X�[� ��)��~�Yq��� H�(݋��{-����Y�t̗�7�NH��Ȫz���B8�g���Bη����SH���`�6`=um�u��
�O�dZ� �z+��~
��7o�O-ݲT�����}v9����Gc�����:E�>�o	8w��L�HK��>V|"��K������*3f6V��-�o���ξ�h}�����}�*��!� ��a��~}{L�� �GL�RZ��^g� 3@�#<~Dc��LP�R+��� @-���0�+X�MiG��21AHցQR�̹���wD�ĠR�~���cwm�U��nV\Kl�l��b�v&��a@C/
K��k>�y�w,9� ���J�$�4�+s�Y���dډ8��59s� ^�b���,�3ĉ��kk6��]uy�9�X?��_��"gL�#��y�&Ͽ;����d�Ae�z(,�[r�P�-U����z�`�樬)רf�+����$'�κ���Av[�b�ms���N�Zq�t:1l|0j�Z��^ \k��O�!'�_����"���:�?)z���L�7T�S!ZH�z?�t�00r������� DO1O�3k��n���"�t�O��O���V��C���{_��`�8��M��X1H 6�6~y`N|�^Fez_O�^l&�\�p��i�Wm�J!��m*h�8�����iF\���h4^3*��_ߍ*�A{���LX?�̔��=}�
� q�7K�����bv�0��
~{)�_Ȟ5U悑O�7��cN�2�7�aD�G��9��ݯ-� �4���y������e�]�H���I~��O�Qd�ZEI@���1�GLJ���@�e�����(�h�OW���D��� �2k�@�&B.�\���!z�# �ٟ��;��P�u��S�#'��\��W��AI�6~�����it�I���������w�E"�UR߅����!Oo��Et��F��uB�X��j*��\��J;�V'�c#���L������V�;7!�c�B6���}sk�b�]HD���o�d��9 �ց���L%+�뒆����'c����cie�8x���ӆ���}��\��� :��7�gd%�2�
����j\���'ϵ��$`I��;Xs}ٹT��%��O%�亁��wg��������A���q�J]�p�"A[ �A}�!`<�p���iR�������޹���A����bW�dJ}�5�u��;�S��Kc�%��GޕS�iU<r�J�?uj;��*���b�6l�=u���_M��B�\��c]aݝ6*������":�!��g�ҹ�=�]T0��,��v�Q��1��owWpP�P�Y-�����,�f�fV�5�I�wK8�.����G@K>��R��IF|י�C�[�
��\��'��YՀ=$cvO,��L@E�  ��᳇�n;,��� �4���n��Z����lO�P�����K2$�p��
���b��*��#��Υ�.Wl��}ᖡ>��ՍNz����W�2L�K�)b|�z��慘���vv�H\Sb8�5�1���p
�8��i%��q'y���ۼ_�h8���6�b�hм��s�"�V:5Uj�"�4p���&v)����C���=B��_b��{}4M�id�q�s$(��>O�C���+L��%&3�%|�e����VdP� ����1��*NQ}�v'�^��!J�����\��g`fȑ՜����6n���b1T&ދ0d,{�
Թ4�lP҅�.��l��"����#���ҖB���Әaaag5=�[���eD$�'�'��f[,�x��GV]��T];���\�U�*���̍�o�d�,H[Z���A�Xfʖ��N��B�K�m+�_��B�OZ2��s��C�C �'��p>ۄPc��sL��T����~�dq��2�|@Q��,�j��Ell�X���0��/6f���U�������P �D�y��-3�Y�%AP��ߎ�p(��'�(��|dq�%#��;l>��K>�1��;d��z1-:��
����O�_Qf�i��s,���Q�m��ZJY�+<Z9������i������M'T��;�s�\����2g�Ðl� �iV�5�qsC3��K���01}F�4wd���1ְG��m�����ݡA�2�����.����Yv+�L^��v�+��u|�|3��4��������,��'�c�.B�cNN� z
�d����-W�yu���f��<}&����X?�y����4wH��C�`�ɯw�G����=uK�Ф�#d��ξz�:^��O���w��;�lh�km8�/����ɧ���NI��V�|�~k�#��v������k�k�[-I7"uf*	��� v�i�Քk ���(�0f��"#F�E:P�;��1S9�&2�&�5s����D7?C������?���K���
w/�3Xu����x�����2���R��	�-e��7,֢Ʒ+�ꆓ��6[aF�����+b��鰂J'�/�ފ��a'u5qIZ��@�̠���q�[��wb/^1����t��6�M�^5�%~�k�dx�r�Ə�ۻQnvc�׌�*�S�S}���,0Bw:|���m
nmun��# �,�F4<N����#�t�J�ף���L�ۈ���gaЙޣ�?Agi�D$s���Rz����q��:��7�|n퍰כ���Ż�d���:�UOQ�����w��lR=&z8��l�܈Q9,q�Ĉ�q;J��>��m��%D�?�G����+�����Q���p~���/)�#zO�]�֭<
�����]�F�Q��,[��,�Tq����|�.m*�xP�)���,H�vd���TG[��$��	��Z�l����@��X�d�*5�7Qs���lߋ����9n�ߝ4�N��>j�ǘ��d���Ԭ��b�w09��>������Qh.}� ?v���u�i��v�����B@���Q�P%`��!i�|��.��̺E,�݃-��j�wⷒ�򉵸���ԼB�����9^Py�޼?�U-ZX	T�P&�T!�N�^�)��Tˮ�A�Ol0�T�b'>�sV=���(����m� �}��K3Lw�e�y&z���t�;��p����@S�u�ĩ,ư�S<y5e{P��A�V-^�Z�3�:�4�w-z�f���	��񕋛r��*ԗ�j }-�\�g�e�LӚs;˖D�D
����V��~�8�6��C��7t�At�
'��twI�}`�/7�{�n/z#e�$�?߂r]>Yr��k���wƕWI'�":�w�,<O�u���T�7����jt� ����1���L�1u�a0I��t"jȞ�z�v]�G�'���kOaQ���N��§�#_Y�r�4���w�px��l/�Jx�\I� v���F-�m���L���Uj@�#'�<�A�T���1LF��j�����ǋ������v�iB���#����P��˙� G5Jr�"�R��U^d��rH��� ��6e���q,�#�����g�
����a%��� 4�G��Y4VB�C�4���Mipa�ފ�<�)�#%���� ��߸)���W�a������v���D�N�����mR�ګn��w@��:"̃���N�4s�&��c�k\D٥L	l�}�6Fضu����S�v�˪.��*Y�MV4X���*�����S�K�4*zq�;��p{���ey�*31�?�F15�7�R�lq%�$K��-	���%k�7�1��qۛ����v~�C<�&�� 491�zH���w��P�tY��<j�4}ͥ����@�����ƅ�X�òي��MfN�4��{TCRʄ�1��s���#ޑ�Z��2A�Yq&��b|*�U9��<��U[45���mȏˋer����.�]T�K�?�L� ������9��V���8�/�,�	m�[�2��&@�0��(���D��wo�CH@���;D�A����DP�1CCC�|+N_&D�K��Cٵ�R{}�j&��*Ċ������7���4�빎��@�,���cy^)�X��R�Ae	YV�Y�3��k���!y)�V͹�$�^1�Ke����[������b��mj�/�aV��5{P���]k��|��0$W�J��E�!��>�z��k?3����F@�F�q�EP���#��eX�w ��� 
a��������s{��أ6{Y&��7�i�Ib��,�)�dj�{|�E=|{AW�mC�/�i~g4�ހ�$��sT��!Ll��t�0�v�rM9:����+��;�sO����"�rӆ�3? u�Е�uJu��%fi1%�j\��a�S(~��D{�kJ�VS���9���G���Z�c�j�_���~٘��`��Z� B�hW��E@a]	:�D2T(�g���By���Gl/1�p���r�H�z���쾹��-HB�5U<8�37�"fޙW�ϥa�ೋ�������@|��;��A���(�Î�?��^���'�9?�&��p`>�^�h25fef0���sH�ՠ�ܲG���Y��i�|���Rdxx	�x,����9p��k9%����?����_�����-a��=�˜�>�=)�I�%��P\7�Ѡ����X�� � 	z;�}�C<�
ۓ|ZLwwe�M<���X�O.|��O+q��ũ`��:J8hǛaA�ߔ�6��uS%Q쑆��6�_�z������"+�����AF�A`6��UNJMق֏�d�������x'������.�
�R��bʌ@�B^D��0���d�^�i�؅l���ˈv����;H%���Q����L����-������FW掆�]�j��BM1|�Z�)
�<�*��y�*��#�V���!C��y�?׾n�E����{?$�ԡ����DD�C.�<��^HCH`ӌ}�y�g?���}C��Mni��
�t��f+ KN��w�x�Z9�i8�w���(��S�n���Dn��LS�ږq��Em�V�y��c��2:gm}�e�$m��K�s��`N�EC���@�b���{a�M���uV���A=�T?��cWY��lh��Eiv؅⫕�̋�H>�\�/��UJ�m6 Q�2~r%��,l�~��W��nhP���	�a'���r�{�aL�m��'��ux��{K��^��ٗ<a�����-��c
���_�\ȏ��f�]N=r�X�/$��#�A�؊���*AP�G1���a�j"i��'?ipgp,�H�cw="�
M{2*��"<)�������X�"�� �i�:e|����D�:�E��zw'�bM�g��x���eQy� (�����@��ׅ�4��7�����OIK&�~捌�f�Ʈ �^����S�l�;Bn/K?A5F���'�_I��p�eԪ�j��}�7�?�o7 ����L�*��3#�wlR0��荒��e��,�������ށ�n?�HI�_�)cH��6������j���Yă[��-��2�	GP���i���9?���6K��J��I�0l���������{��Ia*?�0>�J�{\C�Z=
�,�cڇz5&j�ė�4g�,u�QOb'-!H���a�n�$�x)��m�ay@gT��$��$�쟸�����:��z�I�Di@�~�ϓ�=>���r��_����2�W�#'�@W�GvY{�-~����,.�~�d\C���VC�Y4o�o�R ������Τ�Ra����u+�i�:��?��ڭ���m����Yf&B��W�k��v��D
@v�Z�#��Vu�G��ߋ5���$���R���C�-r[W��v��q���HF�{l���W�q�Eԯ�`p��^�IĐ�x���m�����2�k=Mn�먟�.#˲(��y�o�{�Z)1����Y�=�q�Y�J��+
[�n>��K��6�<?�k��,&aЬKOL.��0��}����U3��:\Y_�Sy�{k����!���md�m��G�͹�=����h����;�
� �����Og���f����w%��3�K3&w��*�m/f1��IA��Ԧ��T�aH��[ W�޽�Z�CT���fÜ�X`p��Aj��D��BwL3�{���o������l}�̚_�?.L�f��{��J�쌎}0�8VWh�V�Y�����v� '%9��I`���K�oy�VOV�s��6��'g��&�IF����փJ-����=E�8�9�R)m\����P���ɟw��FD����p�?� �)�U��-�h���㕶�r|�:ë5��g
�/�N$�U3!
�&qQn\={]����y�
���u8�R(V�0�C<��w�R6��#>3�sB�m	�R~���V�B�C�6u|ȿg�"@��R��0���l'l�gɭQmr����w�l�3ƆΧf� ��_Hl�S嫠��3)��"�:J� n2����r"�昤��L}����i�\�D�TS��ߴaj56��a� h���%}�C9B�� -OeY�ԟ�A�ͳ��y\͔�I�@�1MR�'�]M��āp]}�t����o �w��Ob��"k4b����i�R�����G;�(<-W�6��ob�xږ�П�4J��ݐ�� <�f1��Q���'���6��-�&�SE�>ќQ�����EV��i�y�]@��⧆Q�;^��uП��.�揟�"��fF��=-�D�VH��hX�7K�š	8��zB=_&̨ZU�￟���w�xV��w��D/�= ���>(�l�b��­�{�O��~�.
��!g��E'�=��)uHNS�r/`���E{d�.7�KZ<�I-s��,�2�Y.������.ߓͽ�B�s�t)
Z�s�@K�>���:���E$�2o���e�̩��>`�ecFX�^"���[����0+�Qh�ۈ ��������;�
Ʌ}�
K�� �,������)'�<�R�K%�>�oɥ`���g���G��}@�s-�Kܷ�w�N�>O��jN�NB���7��z.CӯAV��2���)�������?��(�mOyQ<@S,�*@vL �Gk���*�)�>D?D���,3W,�`~N�yԜO�� iHOِ�i�~җc��
�Ke'�hm�g�יۡ���s\#��B��@,\~��x��P�"�RF�%]ٞ�í~y�6�Q���Y^���R�"e7�Zu<t�4�l��:G�P�O��Q�j��L�B��4sWdk������i+
ڋ��������jpQ	Բ
�(P�]J�����{Kr�`=�c��j���e��2�I�^��`k�xX�H�M��6-�34V�����]`�]��6e��`b���0eQz�{\)
��@x���G?�b�t�侒�R�.��lpR��v���Ť%��^���Ŧ� �-i)w�i�l�Ag�\;�|'��dJ��<��/�Ȃ:�cײ��.�/zʑ�5�&X�[g�	����©�| 34�7A�͠T{P�R����$�2ny�é�'KT�g+e�2HKs?u9n:���܁��g؟����ԛP��`��k����O�竘0��z�����j���H�������7٩K��@hf9D�1o��k!�.���||Q��k⽌���o�_��i�F��$�I�U�Ӧ;;{G���_sB/�6���mm��p��;�h��ИqS8؜+c&���r㜰����������F��Eb ٰ�.��s�����D=�+Pa���M�TvU�A^�Vc�"(�-h���9�vY���J�!�j\�D��(��Y)>.,�mE]����T�|�}�x,(Q��,�j��)�b#�GZ��oX`P+�jD�{h����_��cv�@d���o6Aϟ[����g���f����a�p)X���z�§r�y�����	��
w��p��Q���&1y) �\��
u����0��V����/ƐtM�U��'�T���׿;�[E_lC4
�v@V쓓a7dT{O-�u�o��E28 ɮ�p�~��e��zo+��J&ո_�}1�g�YUf5�Q֞�](���%������������'m�#'�Ǹ
Y@v:8U,�7��U3 �H.i�1n�5�v�5l-~}={,a�z�����R�����Q�c伷��-'�|N}����MZ��'M���G�[،``f����=�XlH�h"]�EA	�r y��� =8s�H'U��uS��=Bx�@�cD��֭|�Ka��j�=�P�8$����B���.ֹ��a�9�b{W�n�^s��a+��X���$U%��0���묁Lj3V���57���9�p��bhu�σ���Y;.�z��5��8�N39�v�Ȫ{ch��w|�wi~�W �Ih�'hBO�'���H�ss����^S�u��-~�/"La{ޘ�BcJf�ޛ�
 ��z�Vq!�|��w?-@��P�d���RFm(aP��p
%�ӱP��D!�;;]M�F��٦C�.�o��@�f0�ڀR����Kɛ�W���t��'�4��P�$�,
�A��h�P�.�9;��dtT1(��YWl�T����|6��8s[�R`Ko��4�������L���8�6+s��3P^���ӣ>≴K4u�&��U�1>��/��D�H�GTp�lM��/
{�VA���ޒ�U�[�-3���dm�U3������)���M�����os(�#:�F� :%*�Ys����ڥH�`�RI]m����3%�Ҩ�3L�+A��T!�2�*� 2�?�V�J^3�{�e���y��/�j�O�>9#���'|�(��g��w�VGZ��-q��_��wLGYO�!�6'��ˡ�|�w6
$;�&�Ӄ=���Q��k@��1O����E�ݑ!��22���ʫm�,~�jc-�o�X�KN��9�H����!z�o��=җߞ��=C��P�ʔ@���i1U�ɀ5��7g�����A1H2�YNG��(���ۑ�x̆%S0c�!���2���O'M �t�B���Zx������v|�b��g4���C]�᠁�?ÜmܮxM��ӝj�(�|�{ҕ�z�4��I����Yg=�eۦ��E_&*K�w̿���7���K,�k)�P��j��\�E��ف� ��^*ˈڂG#G!� |?@�(��$ҷIT�|ʕthD�)���f�-����(Ҩ5=�R:8W/���-!6KCixQߎ���\��Ï�N���X�T�iSQ�햤C4Gʫ�c\!s��{iW��5p���	�ϧ@����`�#T��ܞ�X��f��Р�'���[X1ۏH�'����*�$\Y�T�K2Z���6�����Q+I7R�&�,?^�e��h�G���r�0�M�ԛ��-/(�x ���L����e���M�#E����x	K7~�ӔF�� �pJ���/k���l�Bn|[���͝wMli�:��_�4��<	Ơ�,3�� ��!PGb�B�d���hq����l9����y{6�be��é΄9˲�y(l)u}�`�$��z�ѻ=4蜽6l��_�ǵ����Tuj�:�φ����q};ŭ`p����f[p�MQF�˄�p������U����N���#��o�Q�㝉i�`D]&~���V��Ԫ��V����狆��<�S��8W�?z<��GʠQ?�}٨�o�8��7��W��E5a����>@�<����ui�)�^�' ��8>t�͡9�u��<�J\/����p5�~Z6����k����f��3z�?G��~�`Fb�J��K\��~q�B�_{G�|��e�-�Pcr��R�(� ��q��|�7�L�r |���uX�����V��[-�$k�v�u3��h�P?��?����˺#.<(0q�N��OU�=�ڮ�Ye�V��Q7�]e��䷖ʵ}��%@-z�q�A��5�cS����s|K�un����>k�?�F%�\^]��Wp���[Z�����d�+�f
�ft�B�ʁ�*�jG��la W�"�3�w�UU.w�Or=n�j����F��X�ժp���������M�u�<8$̦kH��t��ǚ��bx��$9�w֣�wD�m��Z3���H	z����}�Id��9{�$	�Q��
�`�����e_�Dڰ��z��tS�$d����`� 鬮�'����������S��3<]��yd9�*�K��8.vl�Tj��k T�V ��������h1+���C���ue�%��������QC~A�DE���DE��`T$f�k9)��,����\罃�B��B�:�[ڔ+4��^ ;˶H�-�9��]s%�B���L�ù��\C�����	�+���Ǐ��<�(d��Xg�g;�pv�]mt��r���Mְ��©��$�!��R��Π��������Da_��;�}5������
�����/�~�l�k�z��?���?g����w�Ի�S7U��7aS������x�W�c:��i�������p4�C�z��f/%�6/'���nM�*������J��fN�t	��D<�-	q��j�f�9ak�����Eŧ]���>\��b�M�QA�&P�S�r��U�$��j����K��<@����/��(fL��~�}�C��AXX"�X>ˤ�d&��8�W�R��+%W:y1�IH'�1�H�J��^���MBD�J)k�XR�3]dV�Z�`��Uԋ<�ǹ��f��VI{�F.z�����Z��]aE@q���Ҋ�lUg>��ڪ�v1���߽�����Ү��<��I~;��{)�%O�j�fx'_ۗ����b�#f������9�֯9�r�[[�����+�A/�Yl�ˤ3�����'H�u =�D�����~��bM�.���f4'�IQ�L	�g6\��#1�S1�h+��$(�CT'���o��֠D�s�����|V�x?�96a.܊a��gyLE���R����]l &V�o9�M��) t���-*�7mH�=��O�	4�dl�X�d�L�������B�d���i�jp��"�q3�B�+"�����i�aD(>���ǂ�(+PT"C�����lw�<���2���qh.��X�69C8T�1ڇP���n��u��c�,�?� �xqn�9 PT�PnĈ��fU�X�U�������M�A�_{���YN�t�N���^>7�-/b�KX�����6��z��W@��;����������� ��a��U��c_٦�� ��&P>އ�������ozu~=�5m���Bцbցr��E�
U"�6����m�i"X#������x
q�FN�-�F��s��m�M�6�w�g�!�"����Ʉ�n�E7�
�D���$9܆	��Đ�g�6�\xS\BbQ�@��q#�f�@W�$lj�g�ࠂ�U��Q�YTh��m���PW�9�a�!��7��O�<|���q�Q��x��}�N$�^�q���IaT~(o���#��D�q5�8�p][��1F��^t��n��A�C���PG50fp񱛍hX��F�圾{l��Ů�es�3jiuHODa��� 6H�\�_$�GŦM�b�4���Sp7���.�� ��G;��KSa}�^��BR��}�����s|��`ߺ0�wa�"Hr���y�a�ɋ**j�7�1������.Z႕���aܓSHe���c̟�#�É���Z��H�C��h���H�1FR�k���s�?iQ|�o*
���zfEh�P���T
 ��<ۈWmQ�<]@��.���I�c7S��(#J��6�}������i�Գ�y(�g�:o�{�)p���d6�����C����P)]�"���i�a�L̾��㭈�Qd��ê�e�'{���s��R��Q\̬|�c׈��C%.��(Z����\^wNcB��Ƙ5?#B:�H����� ĩS]�2T�X�zٰ˼��y�����*�V�_}��6��{$�G��t���/�r� �{�����Td[�&@�?���\��}p�#�� ����J����ϭ̘)�1� ��OV,�� (m��J�Or�L����D��+V2���d���_v�N��h��)��S�h�Ͽ�^�����ڠ�Y?�^���X�H(>�8���S��!+Q�e�ȕŰ:te�(2Į%?��i���+L�i�.������b�^���Rj˯%5�SiL�F��]�ʾ��m T�ڈr���eԒ��i=#m9>(�o��MF�l59��p�l�����
X��V&L�����B�D���o��
E�A0���-4�l�S���Y̘x]U��=%x�U�C��8�ϒR>:�DWhh#^V��H��ǔ��ɡ���^rC���Kb��4�Ku�شFC���n��R���0H�n�����7���]7Ģ��^.ޠwk��~Z3f�:(����pm����ʪm4��Avr��5�pk�`��PrJ�ǟʧ�W�gc�H�A�蜏�>�>+�'��^�2#���U���Aq���3���I��+�6Q�ٵV�C-����D��1=wϛ���n`p�TOn���u�������1V��D�8����{!F��8{���B�s��隵�^ _�i��B݌�2һ�a6�@��*���m,�b6�S8�#�jp) ��z������� �yl�H|Wl�(�:�<d�ɸ�:~��-��;[H�|$ϩ;Q�x0�Lυ��hG���6S�k�q�������/R�q\tPV��*�z��28���|�n���<B�b��rN��V�y/HL��wk.��q���4O(Q=��x_P6:�X����Ӝ����H���e{E��"�M3�
����:�K=�bfno��n�(S�d�	������M*<�=,�cOZ��{�q��,PV�=X/ނ2E�j���-��[�B�!X�u������un������xٟtG�N��n1���>�j�7�V�nx���ћV��N|��p+:�dv��4�ʎ�g6l�⒌V!�������.z��(��.�#��6I��x�l�qF������;T�y 0l����c*���0��v#���J$&�������t�#F�Z�b8�{��Fe� �@k����Y�I���B����a����-��)q�jx�M}�@k�݄o��������:���{��������d��^��{���Jj���)*~(��7��D-D�?���㢡|�������]?�PG��女�������2g�aj��\�=��eLd�LR��3�Ѭ"�.sr��iи�9�Q�}DO71������>x��5����uD$�a���ڿΩ��]���t*���n�/;ipuo�M�w�(��}O��/x�1�p���
�Xǥ���.ݦ{�"y�����[�%�t�A*��������A�d//��m^	�I��Ct����,��f�OF$�Vv �C�/V�cVgp��D��z1���he�)�HM�+��e!dݍs�0|}2k�n��A(�&������8^gJ��y`�z���пB}��h��\�A���ޭ^�[���ˈV)���0����d��JEQ�5��t5����\���1����c��5͞܂u��S�N�{?�c���RX/΄+�Cr��l*촅CWU�Ё~=��ģH�p�^�= ߝw\,u0~�c7�����\lt	X�a��?Ӧ+e;rM/����}���"�:#���������(^E�K����,{V�o����b��Du�]�0G�:`Z��B��5.���g�<6L���&��_���ȁ�\@���	L��L��������yz����/��4�g����$����TC��ዒ�ɭ�	Dco8y�Sp9$J�0b�jcG�����g��*z�T�0�P�iN#��q�e������������L�w9�A��g �8"|[���
�CX��w�_�J��S�g��P5�,�G���B�[�M��[O��?P�ɛ�Ma	��M9#8/%k�Tr��k�����1DhM��(1<	mEY���$�507%a�v�Ys�C��M��㤌Kھ��ڟ��+e{�#p{QW��Ɣ�T�z�^ygT{S��Ӷ��1��E
���5�����2�dp���}9$D���C~w��9%�5�Ԧ�����3�Ύ�����4"�B-q$��14yX�q]�Oےذ�[Mvf}"M�"�!���� ��:?&''j�ܧe��9P�Ϫ���߻�O�K�$�=<�#�Nw�gȊ܃.��4����z�,����i��z��O���\�NW�L����/H�|�ȃ-����wz�D^nhw�����k��/��t!6�ކ�X�����������~o+}?���My��,����3�>� �6)FV��G�;�nf��@ UDut��毰|�!���u�@fc�(����ͣ?ג5��W`�V�����g�ѱ�U���J�,���ȧ���� ��!�*|[](L��r�rN�NK�y��dg�L��,l�̯�̬��ǂ��p��T����Y=��'��T�Ŧ��w�C
^�6��^��̭ Z �35y��Ȫ�FrE��y��.ǉW��V��B���Mo'5����R�%�v0��V�ݦ�������t��I�½W�y24^����,��@�~�6�~���ͦ�=�V�7���=���;I{�>�ݴ.�'C�R{�1�D)y�ׂ��kV�tӸ�Vv��A��S�UU꽖vm�{�n�Y�X���1�iS�ox�#,���SP���F����ߺ�O�w��Ȧv.�lH(�|BF���'�^凓x}����iɧ����L
�΃������_��/d��Ӫ 0�3gQ�_���1���DsS��B��0���%tW�Yb��AK&���K���@� ,�kJ�(�[�ᛰڹ��ɫ�\4���7����6�=f����R���G8%X�ʂI԰ �Hr-�o2��7R�._{�I�HJ�� <c�e'k��27|�3
1�zj����AdSo�r�OTN��3B`��[��d6�R߷jT�1��#Q�� ��$<�?�x�Y�Z����8�@��KA��2�u?��/���^�gWy���ʪ^>	�/�f��V��#U�[��pts_?�l]�����Q;k�kq��B����2Q�ퟯ~�L	�/Ȩ���]fXi���Ws_����|S��0V���H&H3��Ux�BC�ʒ ��o�Z�[�������AQ�x1�o<��ݶ� 5��3�V����~_�R&�G)��+=	N-z��%��(�,��G
�Pst�o�gU#��P��0��\T:b%��r4*�<iYϛ��눨�=u�Ih��lFE�T�[�^��惡������\Y�aB����2�����.G�2FNC�u	_�"*t����(�+S*��/��os7j;sʇ����n(Շ�Z���B?w�?�
�qs�l}��/�>�T��1Z�[6g��Rf�=�x81��4������s�D`�Ѧ9���4�tʖת�	��D�͡�Q�d���iu�LG�����<�nW��lK`)E���QP������/�S��gVo����;驝�/NGb���0@�5��Fa ����y��.([�<� =���e��No<��?(~s��
����x�enF=�1*9��3�h�;7/�Sv�K�DI|ö���=�F��f����
��mUfK�;��T�_�u��,�%�^~��Ж&��6����xq�w��9fmmĶ)I�9����Wp�.�������$}�͆�V�x<.���+�_iBY��fl}��|�n�$�6�C��[�:,\��g��#%���tq(����}��GIL_eсz�I���
^����'P�@����ye�3^�Z��]b(ο;����^�|�z��g��܇�1߬��1�WD��w5�\)��Uz��w����T�-f�-Rh������� ���Z<%�H��N�e�q����/��y{a�}?�Y�Ӭ�@�c�z֒��j�c/�h)~��Q�P81*����n�1f�ʈ�K��F���yz�:�h���g՘"C��i<Yzr��?��CN��+l���6G3=��f?�q�O�����+8�?�O�"��r�Cy�G�,Z\�{��gź|\yUWeƫ���Q#��g�	���m_-pY�B��v�|Ţ/�z�!����Md.�^Z�c���7�𰥠|�Zם�0�_F/% ���n�SN����a{����:��l����h�v�l�7�>r.e�ˢ:�
G�:���cU����eޞլ�v[T�g��7���NM1�mT�zT/��G�	9�@�z�܅��X�e��u������)�2E�h3&!��D6�.�7��-��7��EC�5@��tn �K#V�� <F\(��c�	c�E����il6H�~p��S���KJ]�q���qϢ��ƶ� 2z�=��ׇ��V�V"��P�d	��껍'��,?��z=K��v�8�~f�v�T�K��O���.�]w"^S7B�.�_��.:�ѝ��og,6|�hd���h��m��=�U|�ʧ	Zk��u���VL���Dͅ��blX���� z&��2}rA��;G�g�bhg�qh�U�s���d6����0���?�e��ܛ[�?���������k̇#���
Ç��>޳�o�P<NfH����r �X�� �Q�^�����2^�n..F���Ӓ'�Cƙp& $��x�ԁC��нcTQ(�d`����LZT����u�4	���I��&0�l&�Sp;k7M�5K�@GC�h��X����j7Ky�+��=a�l�	[�)��2V����s�c���L�r���}�5��p`��y�����c��6|]SU��?��h<X%[=ct�pC3�н$����`�����4C?�Y] ��)�Q�R>
Ԝ�����JZi>T�-y !���(�����s'��>�V&�� �t�2���4�3��J_�5'�[��l����2�2���N4C�2�|@�$���m�~u��� ��8P@A'Y�Y�����оd�m����+Q�.�J梮?�(�`,Tv4��*xU�1_T�c�O����Ha5I�<]�v���a 9��Y�Ҙ�k{�$~�߱�u	��Fhɂg|1_Q�������8��|ӣj�E�=:8�J��K��AX���A�G��X��4rס�1��Y�ὃӀ�A@��Y��k��� ���|/�9�͟�@Y�ӎ�{$G�~��I.7L�v�|������.cO�Zb*��f_1\q������w2�~f.{���nz��U̺W�I��o���&x�ǩ���3\��;l���r����cԁ�(nu'��V�݊�"��Q3 +{�W۵��6ػ�F&�1f4.���/�77�yя�<ܒo8M:���=n@`����H�q�h�hld
 %�H��Dbɝ���BGۄ��k+ �:Ψ9T���"9��� <�����5@5�3b�" ����>���9 ���w���I����y�����#�B� �k@%)�7���1K�ݗ	���g�qy����	�چ�����V��|{�{��Eg�%���6P[� ��S$��w\�r�y�@�Z�R�YO�(ڤ���_9|��Ľ�\��8�lR�B/ʥS�د�~��m.8~�#Խ�L�G�۬?�|��}Tg$�SW��ml�)_A��l�-c$ʖ$��!��C�!��@$��kj�j�I��A
��ڋ���!������>�͛%!].��$�'�τA؞1A�q4m�gDYo���x:SF��e�+��~�)����(�9�w����Hmm)���+2�[��p� ���o��Qa�_��'HQ�!P�{��_��sH��^�gL`�0��,��j�Y%>1��϶���X�M#�\T���F�W)�-�X3Nj�#gap$��H�Á|���$<zD�j�<̻/��{�JLɛی聽�=�⢴>w����/�-b��J":�\ܢbŇ�5���΋��S�qQ�&DI]��f����
�{Jv7�l��DJE\�fENntCp+�`�4��aw��}��6������`�SѢ����l����}%�9i����Yw$����a�&�
�`��<i?���KF�l�l�0y��y�y��H5��n�����g���v�|%oȌ90�$f���G�~�\�;b�J���O���jl`�V`]e�tumz�_��!dMkMY�&�Hn"]?i�=N�m���ŗH�
Q�fo2����B��D�0�ȴy��aN�5	6�F�bP�b�i@��'h��7mL��D��|o&4K<��9_k�y\������HIrX��A����œ=�xc
:�ȮJ��#cE�ݏ2��xT5����I"����5b"ᒣ{�����QֈO��n<�@H���1�־.��[�L:�3�Af�G �͋d��V�>�D:ʣٍ4���6c���_;Ht�Q��YAG���2�,�S�k\N�	{XLE$���Ecv��PN�
CP˦D�2?�(g��F�v�s{=J��OM���p�5i�'rc���A�U	��ՙ�q'�nS�/?~�0i�:S�C�������=u�"�G�Q�?~Csw(���]e�xw�'IW�(���J�Wޛd��O&�L A�CVxDa���b��QT0����Fg73���H	���݄}U}�>Y�;��Im
�h�!���t��u8����}�R������Tn]��I�MvZ���F3p���rٴw�g�O{�2P>_H�#$�sg�Kn��e��"qř
&ezC[Im��h�:sNY<��,���S*�����z
�+LU*d�=�#�����v�ob��@RWr�ZBp0&��0Fc�4n����˸�,�O��%��3�l�������cL��OY=��}E)nfP+|Y3��2@�&^���l�T4AuVܲ}���>T��@�-�=���W��m$�v�����[��TZ������$=����O�����"a�z��H� ��4�%��&�g�Pc�K����q)ͽA)�>~��O����AD%���r9=�anO,�b��jT�╹e���Xq8����1�;ޅ_3�`z���طf"-8��1����p�+r�!ja]ag���J���"	�[w=���+3��dV� 4�x8�Cye����.�0�q����̂�qώ��&�?&�Yq�ݘKo�ZJ��)��t�$%�؎Ȼ�8�;��� Ѡ��80�T��Km	n9�I�F���leԮ.��|Q���=�aI?���zv�O�\gM�>T��.=�<�vb\�uq��<W:�s,xV�`� s��?�#o�`��&�r�б�K��ByÆTƸ%a#�s�����nN�h�����Z,�,B���Y��[;4��
�	�ot�����U���mKؐڽ�|���\�~�=E�qMk�6fj��\lL(����P�M'E%)�2���t(�A(�hX������><��\�!L^E�+(�LD�<t}�-����w��$)��9��k�����e_O�>�k�S�2�Y{.�Ĩ���[_b1*�~?$C�c(��������e�K�<T�W�=� ����òm�5Y8����{��V���Ȟj��X�m����t��{?²�
���1�4�OY�[���7V��J�nF�w����^2�g��k�,+s�
0h;��k��{!�M ���U[X�\$Cy�̐��TAG�V�\U���Q���-�(���bƦ#��rLxF�n��H��u4G��Kw㮦�<��,��(�U�<�ȏ�]�=cvu������PCX��Q.�L�҅��^�;/Q慎ʬ����$YD4i#��IՌ�N[��mY�ǎ�O~ӡ�3��[�J���[�s;b=Zcw��X�!
�;s���`qoQ�]7}���8�c5WF�2&����55yGK̃|~q��$-��ڠ��{����>2��?���0i��/	M��m.��@z�r�m�� Oo�-�<�^�ȵ&F���-�y�1Z$7�C@@+��wٛ��͚&��;,f�1���e�s[��&n�g��B�s�^������6o�9��n�H��q�~�%ـ���-��N̔$�5<+�e�Hݦ�`���8Ơ�+�Ͻ�>	.g/XQ�}��a'��'�]�*��G���@M�k���1ˉay� j��),q=p�G�qRY'����6�3��@�{�(q�!���ϗ�����O�k[�с5y�g�]8����/�	]�����SP�g�<���� M ���FyD?��������>�G��!�v�B�}f�����=<�c6[A!c��X�2(.gZ)���W�W2���:��hY�-��t�vU��w���L�nّj� 9�!Yg�::���mz����^�g�1�U}5�t��^��wA��@��hl�t��(`c<�z����� ��KY,�'�?!	z^��Q�ᐻC��i�#s�l������Dr��hǆjL�����֚b�/���N[4�1a�Q�I!�?Ş�����"����)�t�0>�7o���|���K�C�{/݃�_P�W�f?��}�B��=�6mG�p�8o���mfk�h�_���aV����?�4�^m��^:�4r}$��5z�ơ>׭0YJ�H@&M��A�<R��z�r��bL��V�5K8�0���lu�D���/@�P��J�_.fm�}�	��h��7�_�y6$�a�`'	����
���x���Y����V�.X9��<#�D*u��:�?E�Yy=]~ w��tVf��r���G �����ٻd�*T���H�c�R�9�ְ�j�z#7h��O������U��M�j�ح�������M���v�$�TI}.�t��q|g5�>�-�R:7��6��B=e�vz��k��]!�%��Y��i�+Թ���T��c_P|1�!��]5PT?NK�6!��E�)�䖜�e��>ܧ�z�u��l���)�v�K��S@��<ʤ��Q�߰��^�L�W�{f��`�BuP�PA�Ƨk�̈�kk���9�b�#��{�3^�J�᱅h��E���w����`�wp*Bm���u��>��k eM3,Ks�Z2�0�w$!Eߌ7�E�ܧ��rIBWL�R�v��%�!��)F�<c�;N��
=Zxv�E=��\���������4H�G8���&��V&�9lʶ<��� �%e_AhKq��CG��P��zG�7�� e�A9���'s�J��m��Y;ت�P۷w�ZC��CW��Y�,e�*]@(�����cI
����j������zna�jw��P����C�&�0�W��_N�����&H�"��8���O�>�Xt�Ot�L���?6���3
L������U���8
)�/C48}���"�ߪ"�t�]i�c�t��W��;,�[��VԻ*nU;*�}�c�<
�7���x�ݬ#�Z\OL"�-[���ߑX`�HdЇ�I�^��&JO�t�ˏ��������\����ZG� e�^���c�׿ӁTyX�o��ӊ�L���������l5�`��@���>���Wq���D6ƜkDq�{��+�|#���6;�B~yYAx�1�{-ۿ^_��_i�J�κw.|.<�*�$u�[q��GLDL��5�$,� ��ot�A�%t�[���'�����c}�弴�`>t�1�@'2j%�v:�����w�iX��h��?�ێ�O�y|�8(U�yk�Z�$�n����{fjFN�&,ۖ2�(���i�i��8*��f��m鐼�c�y���\��-qQ�Z#2��{p-���<my��/}d��p��#�)��d��4��*
�
�K�_��Re���s�3?���J��<�/�-F c�ꁇٯa�����8���agk�c��W+N�M�OT�W�ۂ��
��F�H�o�Q��s8�(�O��c�w������4J�����[�R&�Kn��Y�a[o��^����U�gp���*������~nj.fƻՇ��6�2�~1�.��c���ne��3e�8�	��T�d)��G�Oq���2?PK-+�`+5����@�P��SC�/�Z�1a��2U���Q�Va%��\V��,@�XUZ5��2NzP��CE���'$��bΖ� $+e��E��G�"恥i7�[j]�nԥ(�X���T��Z�r�Y���B��Ie�<��S�X�r�)�d�i|1ʚ{hR�f ��,!O�Hz���w�rw%���Ο��\be�&{׽Ϧks���}�g���x��3��u�x��x�K��T��B�D�^C���C6o\��z����Vf2E:__P��w�{�q���4�d��m�����@�7h&|��8�P�xāXU���[G�XS�9/���V�K��|������u;ƃ~�+8}�n!�;��U�dR�="�'����qj[�X��8��h�cѡu������l��$���	��Pr�w%|�H��|<'p*F�ZT��*��+�p��U]%�`<m�,�Vz0�F>!�}	��17N��]Au����#�a�����O��9��k��{����5fCy�Y+�y% ��"�`����qI	#�Ά�~�>S�7o���>��m�)�	z ~�Y�P	ǝ��E�`�e�6�5�Y�z���>��E��ЧM����wP��������^;ΌԆh��e�Lp��>m.+��-n�UQG���]=��j��t�,�Yj�F�G��X�����nw�%��U�aZ(8�����c��G������HLo���8M��X�����/�.a5a��<�kr��K����;$(�f�Aؗ�&���6,F=�:aB+��yy�z�λv�h��q��I�Ӥ��Lp*K��G��$��b�%��� U]�z���Tf0�_#�	��k?�6
\i,~;(�S�F��K^�J:��#S�C
����XGI�ٚPۓʑq��=)ҁ6��Ċ?�4�x&�r
��t���q[�#�%�|�DWv�.Ob�=��v�����A�8��$��>��d J�.s4���xRʥ�T�#��*����"��$\�Ga��8�˳R� ���h3k�K3��o���S��ԚGU� ' �����E�CΒ?��A�7%=���H1�\�=?o��=^�Kw4��F���
��A�g���%
����캝9��r�&��������Ə�GеG�~��$�Ý��k���שv��a�"f�<���Sf�H����M53�9yc��_l�l�ش���v���:ŷ������7&�Gz�V��M�b�}�hJ�Aʬ]G��#���H0dY��}ç�mz�[ͩA�&/��6p"�ȥ����n�\�&@�A��(�%RQ��fWcLZ�+|AwK������R1���*k��.C����s��Ժ�x�g���7	��D����[�Ӭ�5I���O�F�\I���-��V�H���#�9��خ���")cݬ��Z'g(~�Y���������H�#{�?t�٩;|,.!��R�w��@�q�@I�D�@&O��1����ճa�6���:�p��I�������>�"`�u�/�D����>�jn��N���k/57��a���9��b�`����i`x��B ٚ��و��?��%k
|	p��`����D���V��>��8[�5a ۝W9�M��SD�{U1�1'��m��
 )S�O�۶���r�[asS�-�NJ*g\�r�sZ�$/FYb%Z�uaX�@��zu���'�+���ǦVל5�p�"P��Ns�%�o�O0��kO�5iJ�z�W�q�����Ƣ��f�-
�=�����#��~���eu�{I��M���
�Fd�ȗMRbH�i�/��G�e��?��G&?��4�Ayʜ����2�y���	�^Dr�b.t��q��?5����N��2�jԙ��q�K�}6A�<�$���,�ӡ�L���1�N�u��i�τ���Sd�z���5$m>u�����.�kbcԠ�D�)[!����M(��#r�=;U�97�rB��|� ��T	k�59�����h ����Mu��	�$��T����e6��1��I}�S��}��\�����Ø�ǟN�]L�ʸ�x	���7� �!�=�yO޷䭋ߒ���O�aԎT�5Tas*w�K�Z(�f���bw��/��!��,l�dU��?<K���U��Sݮ�!��
�藱}.�J�^�k�d�cA!2\��(�� K뺽җ�;ʠ��l�:7=�G�߫:47G���<i�'7���x�"�<	�%�
h�۝�G��d�Q�Y��X� �>I���tμ�h�V�KL�1�5��BҔpzA�1�9ӝ/<B.c��x����9`��xd���%�X���v�1�R%��اUr�7��6���_×5�hδ�T���a̌��lM��(��n,��PBNRʔi�*�>?1Pi�Tb.7c�A+�p����GA��T�퀒=*��!4�%1�Dk���=�U\����P�M��̓M�����z��^�6k�f��1�x�O��w�]ח����#2ۣu2�[�Hr��wR0�{����R!|ȱ�G0;:�61��]흰I�d�-8!ȪfC�7��O\'��$�x�q��ｐ�ЁD4�Y�J������
�*B���ފô��Ti|�v k���,wd�;k��
gLmz �X��_�_��z�[%:�di�0	U4LL��-B%���!3����^J��wÒהk��7*W.�׋���-<�~�֘L��Z"���"��H2���$u��Ȳ����w�.���%\ڢ����*g��K ]k����=�N*s�
���x���h{8v� �X�2�Mֻ?(�C�j�xW�f�#�dC�XL@�7�V݁�2�a	8|K��#u��h��~i��Y�%��
�!������=����dbF�h�N�f?� �ۈ묷q"Cg�j0X�QIĆ�L]2�>$���!N�@��ASϛ�S7
��##�؈t�e̶h��	ȄC��Ȱ�b���9��bwZs[�d���|����|^ɍ��MJx�O��\�!��p�w��]$��^'ڏm�e��Q�Qj�f�D��4��I[J���7�4�Zph,n�s`�E&�e��j��*��x~h�3�+���
_ٙ�B�#����T�YP1:ٝ'�����X����o�[1D�Ea���)��<AvGm�ӪJ��Y/k�K�ځ��X:p\t5Ѥ5�Q !�$>j�3O0�d�}X�U�&m��Ӓ����lB�Eb@������L��%3ʞ�x��	�>�5�h�%��x����6d/�^�|�nM�A��`�4���B�!��d �C��+���v��d� ^���gI8Cj0��S���
�����:�M�0��l������ײ��[���j���VS�^nߪ��):������U��r��ˆ��Z|�y������{'��.��_-���1��e)��V�i�{���W�B��D�,���C�aۮG�'	{�!}V�������b=9���I�w�	����װ����''����7�3%��Q9�G8�vw|Q��z�t�?+bN�c�[��C]$����ƣ����<��M_%�������^7�A���p��F���Z[��L�TR����	h};i��a��MEgS%5��~��&V  �jн��G����x�4��-1Y�~t��?a�PrNV��#a��K-ۡLOK�{���E���J�ql�����|��.M.-�x��@����p�e50 ��}	2
�^�M1����9������G���r7���z�!��E�����j���+#��9���_��`=�
���`:� E�W\- ��l���E=�´$@�n�G�6���E��/�@'�Lч�Gێ�D�BW(x3z4h�*>Tz2�F mgY3$��G�����"J>��|?�`)D\�������ץ����n63�Ol"�֓��yN�"��\t�#��Ud\p�8.[c�&gjP��Vm��f���@��o�t����W!�EL&|�����`�<����@{�;����G&hO�T���f^�%8e�_��-�;F�6waF�x���CK} u`��Y��I��>��[�����SRd����
W�����)����8li�[4£ER����'{ĖfW����	;
�b_}�W4��a�:�I|��6b��.+�M|yw
=�
6j7�AR�z_F�E>xe-"��9�WTg�f@zN�	hW2��b3$���K��+v���{���v������%�Cs�K)���,d1��xs�2L�Q���C�ۓ�R׹�v����y�~��sJ<�<���E3;���K�
��/��0rc._�7�bxp�$D4����Ɖon��.���X��Xb"�\��U3��/g?�hqˀ�{)/���rlpqW�/W�s��U���'<�"F��vL3���<���}8m�����6Jt�pcI�Ν7�h3�Af��&�÷�y�Z;Ez��S��?��Óy��T��dn��TgF���yh�h���O�b'�Me�W���꿤�nK�z:z-Qbf�h.緌F~��$����j��E�e��2��x�2�A?�~1�0tda��[N	n��<>��]rW�G��U�Ш���O�*Ć��%��_D����y��N¾��JdC?^�K�l���%��̡,�guې!އ-1��<��kT�Y3��B��/އWlI뛾c_�4��
��3��@�S�E���F�|k=����|d	�����<��)�C�&�e�:X���������I�-�W�_p�x��>�9�Z�fo�J������z�ܛ.p���렪�<Ǟ=$�n>�{�7�ϳ7*�x���eá����o���U�5�>�6�|r��7le��� ���^ʼ�M��p�6]��-���^$�W��nn�����(�C�7���������P�!C�P#fpma4w
J������V������@�dC-3��c�^ES�����t9�����"�1H~S��\��:����l�a��$�/�������CM�Y�eq�1�-�Z��b�����1�#"Zh*�]���k���j�4:���v�	��-��c��x����4���5�<&�b�~�� �;>�b���0�w1���ڂ'N@���0ZRZ�=/�&1�F޸�3��%���Z}��u@����y��zlP] �:|:�O���x�;�1��s�x��\�,'�^��������7�lG���@�O�Y�y��.,9�b}+�Z'�m�cH���s�r�΄����a�N9���r�}|��6��+oP��* �^�ˆ����|�K�Y 4�e��!�ћ��A#�a+��c���8"�q��tJ=I�ᆹm��`+p�&>�NȜ;K��<����n8a��෈�Aoygg@�An�%�ϧ�'��?������_o�|��3�G~0.$����+���EG�)��5E:m��I~vqL�K���� \�b�J#^����F6:C���ނ�I�1��K-�f�/!Ru�r 3�.'�͏�]D���B{:T�IB���*���^U{b�{@�N�e6���ۗ�wV	mW_m�����X>�Z�����i�}f�O��9���Fu�|�rrZ�~�;���AW�6.2�s�<7�tp���� gÂ��i���w���8��|�c���|�p��l�q:�S��%��:������YcQ�*l�,kY9"�s���gV����4��9gy2�c�ț���f�Y�ڟ�ʧ����!]�`��� .����R����"��A<	_ �y�U��f-���6���TjI�؊��ŔR���1޵Bt�`��X�D{��9]�`>]���O��Y���ڜyg�3��"6}�[Т�Ҩ�#1�!#�F�)������l�]��q���� a>g� x� I}��?���Ag��9���](,�zd���T��~i���w��t�J�Y)��6���X�U�ﲆ�z��|�V�����&~d�O�9�e�-W��~!����=�n��e4��������`��Pyv��൏��V�9�����\`OA#K]I�+G9��V��"�V9xAM�Գ`�GLGf� =C���#*
�CoN��ǅ%����R� =��gFw�g�8�\ok��g�i�����8�0���\��Z1'���A�M�L��H>ܟ�@U#m,��:����r���o�|�|�;��J�D�s�ú��08*�S�w止Zd��E�X�������^�Y�ޫ���@�ª
e��$����Q Tz�����x�H�R5,o��R�A
z��Z��%.ʝ���j��ݥ�i��9q��a!�x��>I��x�"IWJ�E�!.�Q�N��x��w���G��(Jt =�>�TS�x��q��a&��93��뤫煩M{)v�!�u4��k���_Ч^�� ��Bl�
��ͽ���tdJ״y��s��▽w_u�����w�s�i��{͵��c ��ika�*I�d!+����0:�1�w�aP���<9GG��V�/�!d}5�1��e���ڈC[焖+1�#�K(�Pmi�hĶ�kN 9e�
��z��ש�N�i_� ���/E��<�^�BCm��e���]k�nF�5�_ j9��yg������jW��bm���q�hp���[�$N�^�%�4�ɏZ�w��\k��2�h��%:/8I1YBΪxBuNg�����i���M�a��Y�8]&��˜�ń���ٶ�g�z���Y-V���T�+��q���:Tʭ��`���s�k�y,�IiJr�*�cf�y|�E���H�7p:��CK�x����:��1� ���h?���l�$ �좔�!_�n��K���~btQ_�x\t�����}�"�>+�"��a�'"��)��I95JTLy��KAf'���R��t�(��\� �i|�E�_�����;H�%���v'��:H\ع��.[�K�k�*(�A����˓�{x�qi����
DܦB�-�|��O]3?W��z��0x6�s݆���|o*qn�M绍�`��7�\ptcu�w��x�հf�UJ*	Ye�:�'�C鸳�Fh*�����2*jxS����.��a��A/�Mv�/R�^Feou�,�{����K̄���T�c��|����廜�J��}�/T� Ym�v��V P�ĎE��>$ 1�0|�Վ-�F�h���rYXډ�����id,[��Υ�aǵ���*j �;�v�-�����R�b)�u��)��5&�e�F��2V���h_�"�����d�"j��u3�p�'j�F�.��ϫq,��f��6y��mi���M����N��tXO��gVnvn�q����j{x��f���c�Jt��j�	�&g�w�7��Ҝx���{��� �I����ph/7r=�8�{�IG���v��܀��m��"b��Җ	?2
Ef�Դ���?�RJ�W��n%��
aoIXӱ_���"��E�;�k�b7�t�kp�%\h~B!��#�T`5/�{�D϶pD��r͚�6�2�\�͓�;�C�!�=��� �W|��"�߽�.G�sG"��+/�{\��l�6�Y�@n7=+�Ew�^������z�U�`������k>�9d�.�I{�Jd���%��.
:��,V�g}��a메���͜�Bޤ)9�ynV$�#���E��e#�5j�,��6"i2� S-BυK,:�	PHeӕa�,��pCA�W���\�n���e��[�x�1=��َO��ۡzwb���p��5"��/�ߙ� |f}�5_0���R�f���7���gG�
�'�j{�R��_bJ�q�b'�_�O{�� V4{��1����`�~|R������d�&t�`H`�ox�?�������!&���Q��bLSk�5�.�Wl���u��G�T(�]�\v4p���u��c��u��[fh# �%ҭP+��Z��@������S��R�w��q����_TCh׻L�w�t8���� G�e"O��5A �PeUy��:������|ł3�J@'0SEX�l�!��cS����E������s�r�����0��ʡ���~󨁄/�o�;���u�������,���"��H�K{�F<{^%�� ZT2q����ޟc�@ݬ���;N��P�L����<I�������gI����������+n�OϞ��WE�t`㹔2�x^���y��{���P���B����h�m?�0�$Ux������:_ʖ
K�C+�pv�ӈ�v��Ad��n%�"�[Rn�U�;�eQ����)ɴ��o�3���+��Vp�w���˧�I�uK6��*g�Q�?�sM7r�j��~�yR�-�*D6ovgU�f�Zd���MQ#6��8�H,_��U �X��Bx$V$�6���AW��3�!2n�@��9�_�@,��%Cx��$CǮէR���߷�|o�S�Z �'rL�o▿Tm���-�d�V�J��Ųر����A)E#@'j�����Ǎ�mB���%#�'����IUy梊��&o�r%�˾?��>�tr���{���!�� �V�GA�[w
�b�d�����5 �3�"8H���}z��b�)Fɍ@�����	��5�;fWX#�f�i�V?)���"���?�c�ɒMIoChCl"P����_�}�G�����--3���|\J�J\�Y.�P�b̯e�YM�|�JlrR��w�\\'%*!m*��͂l�B}u cS���@ORtl�B�a�������f�%���Ed�dM=��C� 10'�Vu���7��!;\�?ZUB�Ot�|#�J��#~�������a��}%����Q' ��ǧ7(fM�Y\C��	�����"�;)#�}��N�=�m�r�h0��U�ulWUW7(��aPa;c��	�k�@1�mV���<5�}�I|X6�$@�b�U�<��� Qƈ,eUf�e=����xT��+^J5:�F�GQ��^t~bx�jIZ<�lh�:���d�����71��͉	eu�]X�!�o��|B�q�q�*˚����,D�d��ѪU�Q��bU|�J�����9(j�-W�ľ�A_��Nr�x٥aX����Vd���4*5���"ă[��z3��q��a��b���-�����t�!��{y���b$-E���
YW$QK�Suu��Ӌ2<�9�`h9L���A0��44�_I"�݌r��N��M"-�^o�Շt��sW���H\0(����_Z/2.vh�v���b]��G�58����Mv��ГɛYu��oC��oö}�	��	����t�!L1�.s/�I����#���Ix���e�xyIYA���7�F0$�&���(�p�Z�z��#h�+���d],cx�h�Ef��3:�I#c�� S3�S���<�aF߅p��u\�˼��[<5<'�BE�U�M�lT�jA�vB�E�%��S�������V�d�
.�3���c�Y�q+4�)V~:[���OR�m�k���FmQ��K�7�]�~P�(nF��%��*�+r�T���t>7���}�3#"tP�G��3V���L�0�:,I|��/�'۹VmG9�t�1�sW��h�b'�F�.�H6�i��I�lpf�l2�}��,m�<����+?%,�Z��sƚ� x����c�����<T{)���zh�u��ܻ������!M���z�3הG����w~��E�F�"Lդ��������:,
	 R��M��8�.u���ֳ�*�6s!�G��@�n(����	���N�m�yq;����qQG��@��w<=a��hQ����aҏO}��B E�8ɍ���i������p7�}
�XJf�*��k#d�VE�0<?i�9k;gX��i������Nڕu���sWܐR[J@�>� �#	)+���J`#T�nsr��Z̮�Lv!9��$-��u8q�-`����?�<>8pvp��g��MnyL��/�4uXx�<xSs�j)�����w�y�!�����e�Ǯ������bX��RT+�]���_��`Z���8l;�
�ʆ��^��y����k�D6r#����!�	���n N�)K����%��J!]�(�r���1�%e���A���U�V�7 >�ő��Cy4j� �ݾUCW�P�'���� iKl��@{�o����d�,��N��t�F(c�'�������"����Z8�;8��ؘӯFL� �L\�p'i9xnn�6���O���iN�����R����S����a�i�j��V�K
9M;j����C̊��	�pn�U���%�£j%ęo$a����.�����t��H���k	�����-�p���3Ԥ\
 �`�dd?N�𫳁�^�ލ�tҰ��.�3˂��ti�إ#p���pS��T���@3_����Xij�X��kl'�Vd�N�n�5(�c	�yᛶ�C#��D�����|�ʙ�ʹ�1�f{���L{h�cn��4v�o��Y}�2A��o���R��j_�R��:�56n}k��ç���u|��V�S�����-��ٮĖ����4���0�B�%��k�%m��M�2��#�-=�� &��9��s�Q<H�4�_��C�����ҡ῭�{g�����ZG�\��i��/�U����~�3���%�숧�8�mX�I�'D������3�����#%#�-�8�K�������3/�3��x��;a�=8"�ug~|�o���,ꝺ�RL-b���c|Iz�ᐹREUcoo���n`�E�A���.���$58][xʋsۭ�t8���w	����f��l�x�l>��W�3��Պ�@�ȓ(dk\w o���$�a��XS�/���Ċ�,�t1.��M�2��mO�P�􉷕�j�#22mY��*�CY��a(���:;8r�=jҮ�j������t��Ӑݽ�D����Ğ�����ĲD���6�	�������o���f�mU�P"��a������ �p��v��s��\Qe edw�˷������lj}P9\�����C�~߇2��#���u�3`�� �_��<���7����q]s 	�ԅ +3���0ĝΗL~(�����Cє"6Q~�&��F���(^�N� #��[����!�!���/L�ڽA@�u=�f��r�pu���Ćo�����<{2W�&������H\G3�S��6�l_��xZ�(�GA+�� ����:�1�5�Cf���hx��vd6Aejj�Rd�޷R0�=���Hy���L@�r85��b�S��'7�%���i�"��e���M�B����ˢ��9�Ӟ����<�u�\a!�I+�H�dm�c�:̟G����a���������0/��5m��e�H�<1�R���,�wqw�A$&�?7���W����|pp8���("BE��9C�����Y��V���p�^hܑ�J�;j�k�B�0�3��Q9��;1e_����BQ��]d�ċ�i�{p�����q�x���������xL�#���A����lRh�7���.��,B���}�F�y`Q5b#[G�ޜ��H� JN&�"҄Koڈ�֑4Ѽu{\}�	���-�S�M�:~^�h�K�pX߾��>/��'�*�驥l(�VߍU����S>����(��K�������q��Ɯ��C��2!T�g��!§�m�4V&l�'!8 �@%�ÝB�!�}h�l��0��}�{������0�}I��6����E�ԪGs�`-���FY#��u6�\��t�x�j��>�L������Y��ol��&����biV� 5q3]0�	s��y��q"W�ۊ�D#�*�*�j�-��E|(�ǀB�5�{.X<�&�$-h2x���.I��,�+]��]�V6��SD��F������Qj����kmrlV�'3y��^ |7��-ԩ�v�<T���|�:�cF%�-��=� �@/����f��ԏ�.�9��R/h��MCտ���1���㇕@�Z�ݑF�Xa���1�w�ޥ���F0�@���G�*/����b��=&O%��+h����ڨ]�29@�Pa ���'�J=��'�z��]��%�C�|��XLQ�+j	�҃�3��4U(րW�ˡ�B3��	�n*�U2��^����QFd ,^ ��$VL�~��?8���N�μ�E�0�xG�E�H����ó��9h�,vϺ^Rm�|�1N�U= �%�X!��>y�g��gY4��6g�N�j�k�� ��x�:u�B�#۲�>��>�Z�\��DJG����(D�70����u�>��|��!���>�k��0��T�T��7P�1G�G�k, Ao���:����!��K�v�\��< ^�D���I�Zn���WP�x�(}!"o^�,�Q4/�FH�#� ��èj�7�w!�r�ӷ�����^�d��ۑ���;�����ɥ���K�u�,�γ�[�W!�Y��&�����d=#����G�<���<�:�=��ˍ2��cA0S��CU��E���+ۮqf���f��e�K�8W�'M셆,q6��}rQa�T������\%�F�7(8d�Y���cag�����*r"��=�2��+s���g	��b/���:{NO�xf��b/W�џjϫ�>ޥ��8��ci6�W[S���v�>
�b��Gg����
�@��%�	�xF��Eg�t�����o�K��bA���ϺM�l�IDb�����y�\ΊOg��>=���G����B7�+��?/�p�*����4dY�U&�ۃ��{��ʫ���S�p�c��>�-[����̻H���+/ݛ����^g�X���,�T����n�n��Ԫ�Jvw���o\����P�*�t�SYF)aPNl�ٜ��jn9�"���!=��o	��&��+��ހ-ܲ�z��0�����á�����n��*�o�m)#z�&r���8�Xj��obCz�B���KES�8b�i}��m�j�ۖ'�4�i��-�J��þD��=n��?�Zf�e�)�w�r*]9��Hã�S �U2�)��?}�|��+���~2�􌤱�
3L`hL&���K[���N\T;t����&�o��.`VN��Ā���ݱ�Ɖ�3������U"� �YD7�Az|K��r�yj�G'��Ag�T��dXØ< "6A�4��يX�r�Jij�{��K�����B�z���ȿ�2��G��0MAcI�9���Ň
&��nLN��D��s���uXo�"'��NE�?�0옮��ұ�|�TZ�07M��W:��vV�aI��\h���o+Y��֑Y��=3�;ӐʷQ��$`��h׈Ѩ��=��Ȃ���QO�Q&O:��cCK�343�M#�#|��D���}�@R���v��5qXnY�[%�ћӗ7k}��bY�2X�m-RU(��Գs���_5�/}�^f)2�/q;��bE�Q
��@H3zq�u〄q1��9�	����N �[��j��WyW�H{�Rќ��0�� �3!d��af������Y���J���UGmz�����e��p(���E�����I�X��|�/U@����YFgy�$�TDp1Ɯ�����tM<�o3�RǦ'�d�=��@�C�޿��������P,�D1�c��i7[������fF�Q���Z�΍��tI_��tn�"4�L�l�G=�/��%~썚����=�[u��]�&�( �-�Sdm5a8;�*�OG���H
�	���ho�6�{X^�+Y���|όa�_����#�/nݷ�c��}�06%��[5�jF�OX<�rY��~�QI��+������,!�N���v�|d�|����o{��F��f�K��`�eOj�(,�"�c�E���6Q�_Z�"��M���Kcu'�Cj����j?��G0.)����gPD�|���u�	(�lr^����pǡ��N@d2���cj$���Uƀ�R�L�M�2�U\t��*$��X�ӌ )���Q�����j8@�{��/�K�WZ���B�2�j�ɴ]X��0�u$�\���%�G�}�6MH�XIO�ڒ�e�v��1�`˲<��-<�>x<s/ ��Ҭ� (b3��Ͽ�mR�hz��>�H5y��ߎ=��kR���?���ĳ��X�w�p�"Z��pv�L�d���{W��#�0P�,:q�Z|	Z^}�Tَvԭ7�&x	��������T8�L�T��z��6���ɓ'��h��y�!��"�M�|�y��w3�6�E΄�%��AN�$�y�=�6��­�T�@[T�F5ĄI,J��v}P��cL�+����>��{�(���P|q��+vV�b'K��0��̊�N���S�y$V'E�9iWR2��a�Hު~������݄qz<FFS�f~��U����H?9�،�xQ)K�)e���@'�ݪ5��p�<'���yW�_{���5�xA�c������RZ9,:G�X�V�� �:J?߆�"L:��?�%�Vq��IxD�ݬ��Cp��/�FW݉<V\�=%�H�Z)���	��zp���r���LX����+�<w�^u��?[���9,/�$���n���N�p�I��m�I?�{����e��7��
4��Iп�9Q���9
���>��*ܵ0����-x@�܍Z�f�_T���A�ȕ��%�Q�L�g�y��cB�_'�ܛ�L��θ�� �t0�
�Z���S�E�;^���L}��X6J���^K��,/��Th�볹p�/�"v��(�h۝hr'Tk��=ca\�G��]�+R��Ze5��tU!��A��m��V�
�l~�$�0���1�hI�4�K��3��+�0����,`\�m�u9>ɜ;�g;���<A{�(��jYg��W����OŲ����JwOc���	�L��,�u }�DÅ"���W���M�����m��+��HŠ����Ş�cd�@�!���رO�����d\֍3N�z&�$\)�.�L���c�D{z�biLL,���5�2�Yn��"��)�(Ayl�:X]g �8���q��\EPz&� �!.T0W���m����z�2T�F�^<|���-��L4���!*S���"
Lg*�JA��ju�0������D�R��0����|}�����L�e��������Ե����K8�d�.D�@�����f����{���`#��л!����PK��tD�]o?9SQy����� �A� �����c��|+�g`:Hz���]�K�!��0�����Ti[���Q��	�?�Py�X��19>�a�1(84�6�ІAW��~~��ձ*ҡ���T9�<���ʦ���L��k�]A���V,B����`(�ld����ȩMS8�uy�qg�ޅo<DK��w|a��<���0���m��țw����
/��Oj/�E(2�B�n�2R�*`�_D�KQ#ވ����A��%�-:�s�57����� ���̘ ����5�<�痡@�=5����稽��-M�<��74r� �}؞?]��^��6e	O���?v�-�̌���l�y��Ҍ�����{�� ��r��ܻ-�c�[�d�E]R����e䍖&'M �����Y,�S� 
+��,֣���h�r�KN��t�GN#��B1���_Ʃ\�����b�T+DYL�FK+@h�E�-�ǜ$=�RƱW�a���Ȉ�؍������"!��й̚���y�F\��U%e;��E�x!���@Ut��+�������'��<�=13I�c�\r9k��)��F�4}������%�[E<�������c�n�0��P_�i�R��R�����?デ5�T��.QVq���i���k��\�Q�"S3xU�"��U�a�f��4�G�V��Ԓ�8��p�i��C�L���x�v_e��
��Ƣ�c�k4hr�݊5`�D$�Smh�o�P���!�)�Lϴ�y<�����|Ϙ�[����z�܉_qK�ӽ��n��.a&���)��M^q�T�:����;��V���e�^M���X�! H�yJ���*��9m�?o�W�i�V�HZi8^~5l���
d������V�$ZH'Xhᮠ W��+W�mu�^�]�q
0Yk�9����f�����uhb����T�a�� k���{��4O�L��M�l��1jB�ܗ�O��9�'G5F^�B\c�H�E�=��l��JN��(X����6�n�a���<D��;�ZꞘ�^{� �-��o��ٹC��.�s!�,��Hɕ?Ա���[oP�4U��TCۓ�˜5���lw9����+�Kppd��j�}�?3�,$\$2�KW�6��r���/\~�kͷ�+�X�}"�59gf;���5�Y�Q{���� �7�X{�Ot�\��x����y��ag�$���9=S/���u�T m"L!r�m��]S҅�#�(=^E�X�ؾ.��
]+{���O�M�j�/y�� r<�n'�`۴�Њ�����alb�p���� ����e��q���fPUA�'�i��[��P&%	���+gH߸u��e�ށ���4ߏ﮳5���U�?���a<}i�_�U�EԞ�k��H��)�3o�X�N�k�)�,1}-:�m ��6hiY�/7(�<�;���^��	��	��o�G��B?���J���#?%��HJ�=ަ��!}?H?��r71�b�yL�_޽���P�o$,���O�kތ�k�8�<l# �_ѥ�9e��Of�I�9�Q�� =�K����o�a9`Ś8��J�˦tٯ�/_���/윿ݶ�Z3���9�5A �7�o(K��7=���(->����Vd�u#=v%�c�m�G��
�L�(i�R6�?���J?&u�}�����v�;D$����B[<������C)B�n�^���>ɷ�CҺ6Ԭ�Xݱq+7CU��V���z��ܘ7X���{7�GgK#g?���R������RҖ��	R�z4-�~l���U�j_�\�v�=H�6?}�r�O�x�~F��I��C�! �I�jȚ[���4��H�/���t�?�g�>�V�3=�Tet-���[�A�1�i�4��>&V4t7���>qܚl�d�QC��o��T�J�ס���ԓ6����zw��z?xD~DC�1�p��<[1����"thP���cV@��~��,��j?@�6a~.�P��`��'�V��*P������7�.��JQE����8.��c��%�|Trῶ���E�-�����a�阉+�� j7��L^-�N�̧����͖�9������+��9��ssX�*Ew�C?π�U�#�v���H��ӡ�����3��h��k�Y䌾d<R���g=��,���29��?����k�4cdi�F�ofBI��/a	���n����
�1�� �p�R�γZIjM�q����ԣ���	�+s� �~2:�c":�@!��lང����������킌;ӽ��Rʄ�
��c�q�p2jOb�Ą_8��*L,�A`^�"Ta'���־3��"R-T��|+H-�W�W7�l�t�($��Z�w3�c���4�1m��EjV,���崽�"�i�eO�2fr�����#����ٛ�F���J�t[+`fs�e�����+�'l��D�G�q�kn~bI��P�X��C:K��#��ދ�c�E���qx�������Tm�\��!�Kp�����4}aÎg���@�������}��'W{�Ɣ�
Ӏ�ԪL��A�qUz�A�<g��ոf.qJ��-���4N{��2�P�>�8�cV�Oua-v�U�
��x�%��rg�^�7\B��a�=�x�  Z�թ� �.4�3�:��E��Z�o���g���D�Э\k�v��K�e�}��H7��T���U�W|$���k�19Z�w6�ֿAZ�*����&���*���f��`��T����īЉ��i�%m���鎨�|�ʉj��uF�A�vUؤ����(Y��F�N��	����U��d�ml�U���U������������$��a%�oH~a!�֕x)^<G�$�\�dB�z�T,�K��̑z����'���hu^�G�Gz�B_l:2����`��N2�N{]j�X��?��fZ��-��#�y5Q~����or��@Vƞ��kP�(�}�z
�O�����W�2L*]�%�� � J����7EG��2���!�1P���<�Gn������DG<�L�+��Ͼ�2��=�o���>0�^�ǔ"�~Ƣ���G�#s,=#޶�Q�g<�%��Q�(��z�	~�V�w���θ�����|S%���_��rІ cw�y����� D�� �%�����k9�F�!��p�dEt�:�-*��¹c
��j�Վ�����[�ꢦ`����~sG���
r�xK��Ng���=�K:��Xo�vHv�<���2�b{~9�@�i�Qo��Q����#s���6Is|*�ߨr=�P>�% ee�J��mN�	Y"��򇳞�..)�5h1SP+EHAZXWd"�eg���~���ٌ�r�(��./K�#��τ1J��S}�l��d%�L��ӺĀ�e���0�l���7�S�K��P*c^��lzL�$�C�O�'.*)$�������s�'KmoRX�#I���1���5���q�ﶨ1f+��Y*@�4�����!X�+�.��jGĥ��g��K��y>b�Tь����E2�Ą5��&����A��ꭲN�n�[���T__�.����`(B=�M��L�ɘ5�~�Z�*�MgM�y�͡*�B�
��W^�����{�1������@^�����G�+�|G���_���m{�J�t1-�췉��^ �-��݆δ�Z�U&-2�=��p.�q�H��U��$�Ľ"��%�6�����f���f����M�?\ݿx�����/O�`x�bB�<���;���70J��1q�����9�,��(	;JD�P��a{a�X��s�'2��w|��>n�O=B��z� ��=(��o���F�%����5�w3YH�f+�����������54�^�tgե�m�|R��z E���s�[��XHO��*�g��Ғ�@��A��&���M����� ո!��߁�F=\�*��"��c����pԐ1,Cl�\Y�Ә���ı���5��ɋ�����������r"�k���ZN9K�+�0��A�Wq}7�.�;@{ke�dVF��$���a��~��9m�$��o8t�~�r_��zd;�����zj_$�Pڝ�!���)�,ё��zji��Å�h��Kqx��r{G
O�d�:H���Ҳ��nv�F���dU��]�qk�?�/�6*o4���mO֒���b'�ۍ��P���6')	��v�(�<�����hf�/ʈt�_Gg�J|��(��S��)Uƒ�M��;�9��`s?�*���>��*�U>��>��}��Y�����r9�SBf�UI��R�ڤn���0�f�t.�*��8��]	��#u�_�<9��>�#m1�>u9����=k��uՔ~�
��I�li�Q�6�ʨ��|�,�������A�t��> 3��iB�oS%7E�d��\���aVe&o�8<D����+R�L�-��jX���O�M�9��µ	?�;P������t�JiS~8���|e'y�/8����	v��ta�R�x��(C�'���}{�U0f �nTE��tg�Q� '�D��|�G���,�g��>�ݮg��H$<�T��M6�PO�w��$�����UJ��	�Q��R�H 4�ֈ
�>�8ҲȚ����r�1D$����ާ�ͽ�#���"�)8ɱ�C�ql��:���i�E�gZ<�����X��;���(<�8����з�G\��<L4�Pz��œ:H����8�"�v�ԲOZT }JR_���]&�'q .�R����'���������*��e�!�����K�eFْ%ǼNma�ʙ��*i����p�S�<NbBN�����Ӷ��H�g������W`�;��y��5�܇:dCB�O=�6I�}>��[7a�T��?��Ş{��S��=>�Vy�p}����.CS�����A��#��	=�f���Y=��w8�E�N
�xN��Y9�Pȵ¤���R^jt͇G�2Q�W. �e��nU/Y���(Z=N�-tƥ��w�[ivĹ'�-^�!b<М^�;��<�i�8Np(_bI��WB�7��}���z�g�1hV��P�n�꽲)�]M�����o�z��$�ox��/ZA+GӅЭ����pkG>[��Y jI�OHB0,����=�$�J�)f����k��ᣆ�fε�\���v��(�I������)�U�)'�ҥgN[���P:`�|}[��׶�
����>>?�V��X&ɽ��p��H��~h�FBo,A	f�^���#/@@p$����tz3� �un,���Y�D�)fW��l��N� ����wQ����9���	1ō)�POu���'��y�xLgJ'0U&HP���˥���z��4�:�`�aTb��Y�ε���������h�8�%�̳��0Ho;�fjcT/��Oۦ���٘ztl�0.3�:o`UE#N���W�~�9��t��iX��#��L$�w�nlc��<̐t�TP�*|�6�SF�K�����z����w���y6�<z{z B�gt��Z��F`��o�ҏ3��̉t��[���Y�f�k��tc��',n�#j���L6#ј��[몒7;&}�հ>��;�,�Bb���p"�����>���k��c�`�*On�\L�����,&��16)4��b��NHݽbC�K���(py�Vv̈��0������.��糺y1=du)��� �{=�d(W�1��J�m3��n�ej4m8N�ߌ��=G���"�i��"�f��D�؊6�����L�]m7���d�g��ғD����_�Kx1(Լ-w��N��&.}`��,��� u֗��T[%Y� �"�� �G��%����h,�[
���z>�� ��LB�XrHB2����.�zǆ��_�"v���|��X���.�)v����)�ѻ(l���Ԅ9�����n�k�G�oB��挣�ꅯN:y�W��ٛ�1 Mc�J���OҤ^�:q����C���В_�/g)�BR�2'��D�׍�VrwV����B��%K�� Q��=�&F3B������yQg����c�\m7ڥȧT���a`�e�p�v b�'��nP�R(&�e�銳�٩�f��T,�,����<k���'R��E�lH��>�������s�a~�+��X����a�x��,��6�$�O6�/g����BRT���� Sye`|I�k0�j��մ�4`�ė�HX���]1ξj�ʫ���t�oN��΋�g��Jݝ��]֭�S p݉e�s��B6�l.�4���/; �����1˿����N����!�)B�G�ͨ�IT�s_�/ �čv���6fCO<�?����\S��cq�	o���*\RG7�@���K���5ɰ�,�;cNH�8��``k��J���Ȏ�� �V����+�_�m�r�U�~�O�t��,�V�TN�Rk�,�s��]�x�6M�{�)I�/�wb-��V����b�@e`|o��,�bt�r�fw&�ȁbyo�ۥL6�NT�ȗ�f�R3� _�S�t��3�0�3�/Ob1���@�.�T�Ndl>�5i>�W���Fί쯍K���_P�j��S:��U���cDc&$�Y�����"7� @���u�z�$`�k�$�x��>�DdO����klH�FvBbZ��'��l�q��r�Ҍ�7l�7�Lb��41��Fa� �����+��w������$����	c�0�p�D�ىT�ѫ�O����G�d�"�j���F�!��z��B��R��$������΁�=*;�ÜW93���A���k29��O�������{��:��Ҙ�4QD�M �^��f��!��!3)`�3�ꆨ���c<��b|"Q��L�.ENLLjN�X��0�����Z��o���C��b�K�R� �OE��h:��D��G�SK�g��ϝ1[i��VU�u�l^VFC[�_��������$�i-#�cL����>0�����|5��X����>��a���b�Fw^����~�N����	8d3+������Ǣ�'�-�$����LR��������
,v�@D��	��t��P���?e�vV߿aG	g����wvǂb�.8^'�w;�m���k�Ve�׌l(��(EaF%�lG�x�\�O�϶����8N��}�|e^�A�T��Ib	�-��e�,[��(2͒f�̝�D��D��B
��W_�MP���?��W��5�����7W?�;���$��w^��̞����QB�ޢt�ek�<��:��Y��l*uPI�l[�=/�bl&I�I�>�w��3�"�4����+�����~@?�����^�@�3��������|n�fmiQ4��0z��"Jps���]X�0V��Z�/��s#�[������b ��g�,x�9�9K=5Q�«-�Ls3���Ɏ���(�Y��q���9��J������R�5�1�|;ZȽP�jL@;C@q���wUh�sZ��ј�
���>�f8<�0_l�X�zS)J/ڑE��d�d ������� �x���F6�+*��ּ>1�BB�Um)�%(�|��s���4#������"-�0�x1�Х�_�t��&���k�Q�4��<<�XtA��G4����-��:�$y�����b|<#�I�7sT[Kq�LH*[���7{���07�HC6pL㫨uqngݺ��L�
�U��SZ�
=nTrj�gD44͙�(��^TM��x�M#���g����.�׺�a�L�+ �k��,{,&�1zmk�A����Eh3�IͻVG/+�2����A ���gm/��@ �tă[	����..Xʁ���o�����`���B��ڿ���(����Ʀ�XTp9-�H��k��˳R��ս�{���Uth��g����8<�$�@
".��ݖ2L���fYI��<����"ۊ�t�'_"���z�l����m,H���.��Am�W,�&����P�>I�y�=�>�ږ��ė6��$@I�%
��8uBXeE�� ��ɓ)�]LfVD =Ƅ�i
?hXϪ�����d@�߉3L��"��2�f�t ��Tj�r�?
-!�c*'QN�ão��_�ѐf�y�­{�R;�����R��{D�X�KLNC�HQ��1Pz7��9y���_Dd���-���`z���p���vz�2�X9um��sf݇��?����SO�:��wT��VǤ�����FpR~ѝ�i,�7 ����F�XH/�c?D~1v���b�xu�%_���&����Q?$��ٙ���G�7��fmr9�dea�9`c-7L{yNcy��`K�dS�4VW����y�4)�vMB#Hܞ�
D�W�����[�S�5��{K�dI��%���j��7�pW`g���+�?�0;��[M�hz톀i�O3�٨�"��D�叧o!y�Uf����t�S��{/�����;��xzsGB�`�wԧ7pD�)W�����0���hy���`L�%�twN�\�&�>r��Mn��a��g��L�ӏ�R�=�p��O��[ɽ��u��z8��,I�YGNS�G]�EҜ�o�����`��(!L�Ъ0ݗ��楞�K@��P�76Z+7�Jm��!7�Yz��&zGM}D��K���EL@;�����ڕ�f(������j6�RZ�S���9�i�	Il�m_G"�R��3��?]��*˄7j��]d_j�?�Y���+[}�_[��7䔮m��)xo?_��SΧ��f�jh�P��!��4>+Ϙްs|L�h��%Rm��N��[$�����V����^���7XI1z,�L������r/@�In"�}7^�,"��Q��H�s ]��|.`$$�_��8��r�xU\H�^��8���۸t��&��M�S����3+����B0K�Z��~"��]4��ax�,�^1�GAy�t���5;S?����W����6-�A�Y7˳����2�� �LdH8���UhKi��Qg��s~je��:��7SS-|��p-lmS�ʔ|���������D=9;=�%v�GOI2lsmx��q����>@�D�2��˒�q#h�c$4��,n��+��A���9�l9���s�(�V�
I����[n��
�?��E�c��#���<��my���a����C�uҍ��'AL��[�G�$G⎸[��61D�>�4Mٔ8W	�>�:�e]���gf��ϧ��Fww�]}	�ͨp�Y<%�֣�^?�}3��^N8�H��{o��6*��ߑ�j�=��v�@�D������n!Fz����;��]�eޱ��!�x�bq�N �]`wG?�8���$��m�B�S���g-���aTb'��h]e���� ���6��R�u�.�0j=_��w�3���Cj��8l�CD��PյДCC�42�lN$l�[�|�ÖnI���p�M W &�����)���f*�Ӏ��5|I������f��0<��dws	��~������m�$��z]���91Y��Y�:�	�D��g\t/���y'���r ��B�#�4�bq܆�x�	�?�9�ǔ�-�`|f'_/T# {G���>�(���.�yYx`��m�ߓV(�S�r��M��"��&9KY��P�\%"w�[��N�Pj�����2�/t>@a��Ir���sfT��B/���C�U:
L��
���cy|�
��7���n2v+�����7��h5��\;I��k��1'ד��G�i�0/g���sm�x���tkG$���Ë�f�t�X�h�fD��� ��d��i���A�D����;�@2����4�����-d.�k�H"�������d��	7$6�~D����U��P?0��4 V��Eye7����eɣ����AI���zC�d�
���6Pb�bE*g0@H��Y��9�n��h��kR<xOᦽ�=e�Œҝ��*k��sJ׼�Gz{4P��׋bx���{R1�jAo�3�{I'\l�-��H&~&��n�|$Z�z)���߹�x�.cg�R��c��W�D���`�G)Kn�MF�]�ϲ��ZI�����*�R�	k-v���_F�0O�R����H\b�����8HN�yK�6_�\�K�%5�Z0�S4� VB+���%$���M��3��' I)P��y����\r��'
Eg˄�@��+�z��	"�P�;�G�~��>��c�yL�So�I�& ֦��ɚ����-���>ed�g-gCAT��2����6��G���r�տ��11`�4�XT5�t��BCn��w��f����AJ�i�<�M2� jҎO7{���͡Nn�4m2� �ɽ����b)�k2c^�7�а������ϯy�v������ޔL���	��;(��C�ėME�#���l��^�6R�qX�i�
N�ywK�͏���*:���Y��s)Ւ]�z*m�`L���dĈ��y���䭠/R�Ӷj2��J]�lҫ�E
&[Y!�r.�&�t�N��^�O��\ṇ,���_~��@��1���}8�k��V|���N�Qo7�ʅ�5�h�vc���F��-��[���W�t��z��	Ζ d��kj��T�����Z�c�#,t�kL���"fD��|�y	�5����D�N�b�0]ϧK�"�iS$a�lS��\P��@\���[���S�EB�� ڕ�'����=�sd��v���I����
Y7���W���[R=��1a����d�'�����������'�+��rf@�+��&~�>����Kmg^k�^�(�4_�y:ʛ}���͏_~+���4����r���M�(�ӓP����e*�-gI�D����uf��'���X��Yz��7���B�w�H�,t�hk�e�OS K����N�qiF:�{�vz�y�8�+�&�or&۾T}�\�~�2�w!���D�V�A�аDFh�i�5{�3f�����G�2��㜸7�3�k��}��F���0�v?~ ��g����/���i�sRX�
OFD��R:Ҹ;:Cڊ��DfO�~��x����Ѩ�[�<�n{�/���Her���ݵi��_��lz�h���M�oe�o��k��=n�[C����h�y1,Rb��_T��58O���������Hnv��1\U��%�n�m��S�O`ȴ���kQ�IobR^I;��l�H���F|yǥ��
D� �� a��d����Y����(�P�oY��j�(��4�>B�5��ϖ�Q�jH���T>�4o()�3�7�b�b��؝�|7��4��˘�[�6#Ż	�>��b��2�%9�xZtR��?�{=���:�8����v�f��������̣ђ�X��Ķ��0Z]���%&k2�K���V��C���0G	6,�Ba�=:��S�3�z�@��k�5��Gڎxt��[��ڵ�F�l���4	�E��k�X�}n���<�J/]^bR�	���U_���cZ�1��h���iq㜞�o'��>��e[�p��V���ĸ6��"S=���E�)��+3yM��$�/yI�-XA>@���$A�0D��p�'��!�ҴL"��}�3�Qp�O�c��b�7jϛF���
��j�X�#$S�ck��9�y��9���I���-�Aqb�πT������r�P3����7�6�ٱ��!�F��zc�'�6��^!)�4L3(]�_���� b4�Nn̅M��(N�)��ƪ9��o{�MƇ�ú�:=���q�*���T	Y�v$���;ctӘsY�1# �<X�*]&zy'�)Y �&%�����!A>\GG���!w�8��<�o�s[�II�J?�.�w`Ji׼��X��ɢ���!<꼬C�
8��aH�0��u�D��U�Iʢm:��5pc֏Q�[�.Ѽ	npX���:�T�+:!k��~��4���D�@�]���S�{փκ�����>ٮ	��!8R�]��z��mNO�mC������ڏ��t�9�
u�/���Tm�G)�ר&��ɮ[L�cqIg��%�o���2�&�{4�e���ȕ�eq�����JҡuւȊ��,����-y�p1�;ù�pχ�Y�{����e�"äL�cL�nH�����h��+]�W�I��L�ȩ�'$ӕ&d(�*�L�ִ ���)��_�[�����m���2�<gI�q��Z���c9Ԟ��{�(�����v����1�>/6�����P�#�_�;��ϸ�H�3s$�[�?�f��8}2��E��j\���)Y֞�����΀A��;��^�.оk0熁]�
K��C��HW!��mO�@�Z���� 3��&�jd=���6 ��oU���s����I	&�ٗ~R��&U+Q����CQ!�[
D'�A�e�]�yU�!|0�4�Ԯ�l%wߋ�h��~�(�$����	��Sz�1�/I�b
�����Xt����u����6@��G�>0���jh�sͮ�Z��<m�m=)-��d_�o*�֐�e�#Xfn�eS�7��:���Xx�#~阋n��☧9����J
��'e�!%ʢu���ZZ�񴥂ګ�X"���.��Nxi=�	���ǈ�e��T ��g����=o;�5<�yK�/�!�<h@�ytj�0^T�ncp�!��n`905 k)@��IÖ�^�y�?!�',CD�	��N��)�ߋܹZ��ߠ�m�x{֬�@w2(�h���i���W���}}-�)�j-ՠ�7�$�lN�x/}�)��Z	ǀ�7�<���a���n'�A�hͧ�畈dE�2%�� �Ƞ�ȷD{b�EKD�á��L%�0al_gLK0A�S�ĭ�=luVB(���Î�9k�u�q�	[c�'ڳ�b��R����J�L�)����i���W���.��YG>W���N8!"���R��� �߼��5`�A9�*�RB��-�hݐyTϭh�Ĵ.�b&�8�6�~1�:��)�E�6N++^��8J�t������oAK�����D���`�/PB3�C�>�3�b��7\Hbf@0;��m*��"�`�~a�;ԫS���`C�D�d`���Es�����B�s��0�D.|���1�Ȩ�������t����z{,�K�Kby��~����zᥑ�"+?q&}TeO��r9	�����wya����_�夫$1;��%:~v��i�i��6c��[��3L �m5��:Y! �ˁ,��&�� [��neFE]MG.Uμ�LmW53��a��Ȱ�sq.(�E�%?qk/��顖��ps�ٺk䓰b�ͤ�?��i�L=��
�޸C(���Rkhy zs��N�f�������rI�� �+��ٯ����I������c
?$�h/
6�Q�*�M�����^
 $�	�Dl��'���.>z~J�R&�n1;'�a��ؽ��R� C�ޒ�P1�⥰Hy���"CGy��ݱ��ν?��{�F��&�P�g#y`�us��T�|P�.��^V1A��K-4�������飷���Ր�y=�������� >�y��D���X�A�L2�N����D%kU��4v1��(��A	��"!K!Q�$9:�bV����a�������K��Z;�t�!����i�3v��^Z�1� ����}��1Qϵ�vԛ��fvrv�����V!�h�[C��d��xڀ1 W-wa��l��F�+���!Ы���	3�)l�z4�1���0�h#Ph�+O���v���Y�$���(��,�*���iI��摬��jl�Ƒt#�l����\f��R��t1�{�誄��>>d�2���ELdz2��s��2��VJ|H*���xy^�y�6��p����aZ%�`�ν�[��lD�����'���ߠ��<�	g�A����=���%�D'��M%���9��Y� �:��R�񉤌�GRM��L�&�bb�"6�٧��_�9yF����A{O�N_�셆����<��2B+��g*��^S4�ᘮ�}���-k� ~��3_F �<پgVl56��C��cj�J���| �:w�Jk��L?��K���[=?�ʭR������t�!C�o����W�{������RD�K(-���^)�j�ؖv�9�v���
R��WK��J��]I�L@Q�d��	p ��Y��K}�C�	
�J��i`�N���*#�\�d���ب7�����_��]�H3�#��x��Bj�[>�F;e��$��9��a�uщ�0��ryH�"�B���y�$�n�%]4#WqpǓjD`KR�z	Z<�=^����HY�fQH ����.?��J�������}���eo��M�1��^̡S���q�J��2Kpf>��e@�~aOi�����e�\��I>�����S<mD�w<*X/����N�0y����,����?�}y\j��ʗ��S�ݑ,w���m����ae��l��G�e�����to|kk���«���i��L.~�+���T�Z�� 3��v,��՞/�i!�!�\��#������%	�7ʎU[^;\�-�����Q2
�#k�U����B[����0]ݨ�E�Z���	�S��NG��'mA�	%0G��ž4����8��Ơ�\����4�0�s���:���8aJ�z#骐%ĵ���9�����)c��8����n�u�DWo:Z�Ҧ�le��W\J	ZY�~�������&�uٻZ�V�S�G��y%��P��t����s7�m%+� ��*�M�}�km#.�㣢�4e!�w�J� ����%�M���" �O�pN]����y�)���9O%��8w�cٳ��h=���2�B�,�Y����w��_�:'�k9$�?Ĭ����
V�*'{T�w���R�8I�\a�M���i}�D�`��dg#z�q�z<�9�Mz(����M)� T��9*2���%�b��f�;G��@;���aH(4O2G�=̝we� ��^�謧&�A'~�tQO�f�����(��m�h�R�[�'Z���<R]�0<0"��*��{���e��K���Tx�e\��:���8s��d=�w�����h�  `)fj��
N�dpmr*��NV�wx�rT��d���a��鯟)�@ݙ�7Haͭ���n�����
ŐR邏\�ai�mvӘ����pfg�O74x��~��B��D����z�&ON���q.�]fj�!=�R$�QX�gA��G�aa}n޷0(���䳷dA�`:��E��*GVY��c���)Фw��k�'��A���1P�y��E�c���!��k7j�":��[��M��ߪy�KJ��7ߜ�!'`���R�c���U��q1nǱ�9�#w�o4���l�7eu��Q�����M���ŽS��3�+��9�5�m\*A�3�����8��		�ex�z>�O �e��X'���"�����u�r�O�ك���g�_�kU�x�!����5�9�(d����*-4E�Jt&���J�A�K���:�G�(�H�7vSV��LL,{U�Z��QD�T�ǝ�@3��,�y�@KK��0��E$�+Ķ�%���BH��<֥$H[S�[4�I*`�؄���d<. i18T���.��_r�ph��C�1 ��uڝ�Њ�B;O_��?~\��Ց�1ha9��s��V�i���.xiG"�(֩�z�4O��fz�씽����/n5�ۡ��AZ�9!�f���b�� w�t��^�6 �a�e@��=�T�2��. v�J�?K�����B%&! ;QL��k@�kcy8��RF|`z)�>y�wCR�%�0���d?����||'��L�"K.	���Yь�k����*��F��Kz
�xu��}1��R���dg=X�X�����	ӛ5�`;����,�����'Hmy�1U+��T�~尃d�j�����J�c�Pa���|ѽ�	YsyIA��� ���x�^^�K�y[o��*�r��^l��r���
�������3�+k3���6o���=>y�z�f�XE��X�n.��b���5^��{����w�b/�ɰ	����E�Q�́��+8|��R\6�v�e�~��qL&�Rj��7#�R�A�s��5����Yq�Eb���<K�W5S� >V�j����.�~�eUZ�d=��5]8�"�\�;�*��:�5�ø�d�&y���-����]��A[G�!L^�VF�H���D��`lCgg�<��
���Py_�l��^�,�,��v�à�-�K��= .�*�w-�)}P\i��H�ݰ�B͕���P
mJ�;=�+φS���2�$[Q-e6DۥK�W���^�<�OV&�����y��X=()�JDvہ��8����c{�^��u�T�C�AE§+Ȋ{�/����.�Z��?O�G?�D?�B	|IVz�|È��?U)������[���A8�%���C.:$�	��e4,����δ��83_���p��t�ڸ! ��6}K{�)�F�7�_Y���_��{#��Ӹ��b��B�I�ՃE6���u1f����K��AN��r�w����A"�o��N�ޤ[�����|�Lau����m#�>�:�ͧ�W���o[fI&�8�뤬5������PԱ>V�P��B�vz������^M��Y7�*�������g�ڐ�� �(��?��M�I$iXI��n7c~�{a�v-���5y�Ï��Y� ]���+���&L�$0[�ت�J�n)�84�������42�Qv��Q$6X+e2"Vq�sq11�
,	1x��J�_�nBҍdY�Q���A�~� '�_����������� b�����h����������y��:�Q35]�P?�H��9���v�2KH�U׹:K\Z��M�k��4����K'q} �U*����? �� �7x�?YB�ݽ"�i�����ߕ�xYz�WJ�\u�1�c%�܏I9Q)��'уr֌���d*�N�n�ut	�>rܐ�%��������ȗ(���Ҩ����1"�(/���"��ߤ��]i�"x�|�F�����?�u��r��;j&�ګ� �����v�Z�|�в����$�vc��բI�k]��s[�>������H�/�<�d#���������_�b{U\�<Y&����6w�֎�a�e'���>�F�0 ��#�e�_�:�]l oXB�I�75-��$��y�ǚrY�7��=�~Y��t�IV{��>ı
�ll��u��B���9��k�Go���|�xV���!O�&��=��Sک�ʬ������م��n��W�T�:���#{�Mm�'�S��X��Z�M����E��p�JB�w�[�E?l�י�f�|(��m\ٿ��z�\`�P�)�A��*�����t�X�B��";d\��1��\�F�H"�@>��A����dk���C��2N�R�QR��C@��s�8eH��l�F-�D�x����C�'�P�=w�u���5��M����VR��{:�!e��0�~, 6��am����c���ZTNF��>��xZ���W��/�,���%��U�.����,���U	YV�:�4��7Bt\U�ME���3X��{���2��w���c]?��'F
P����+��Ҋz���+�"��
l�:�F�5���!xy��@���3��\$��2Ow����`�g��̈́��\~����R�&��x�%{��������� �Ȯc���vm��� o�0M*��=���_���s(Pɨ	��8�3��e��O�'���ƙX�u�����Gp�W����>Y�jNKތ21 U����Y'ӱ��!�H�Y�I�R �i�,$Ņ ��\����.�y�ڣ�����.W�4�V���U�z��k6m�n���RX�[ÑBL�9}'��2wm��1l�p�˂�I�]��s	�K�Qx_k3@8�F�`����K�g Q��
ը�3�1�4R���U}1��S7c��[�oԪ~3i�W�nZ\�9?_vG1��_с���d8j,�K���:[A�܇~���������P8���I꼉5)Bqe�Q�w<��`����e������t���%��xQڿ �)ϻ��VR�Q}�﹕W���n�#� �����Se���e���x��.k����Ɂz"�6A7����s'���v^��_FEG�/g��!��0���M֬Λ;j\f��dͷ���]8�NG8D�K���������򝛦'����I�/lfv<��B�ظ�.�������d�C7-�R0�\";<2h#"^��>kɶ�z�yy��-x�U��L��9�!�
u"�Z23B���(�Ò)^4@~�b>e���;��s�G���� F�:�|J.+V@*��ӿ�����BA�1>	�iE_7t
�D���g��#�����H�l.�]w$�A��j�hŲ��L�.��?��[�|�~�~z�),9�<3�N�)5>р�A6e;Q��r.ya����,W�&���0��*��.D�u�KGS~7�L�,����������{��E9�O'�^�_���f�»�4�^ (���9���؄M�M�r���>�9�c�>�����Z�?�lS�٠ǖXж��)v�͈���_� f� �B��t=��kj{O�U�� ��|h�PF�}л�}�@�j��vȿ/�h�NUfP�[�QT+����}�.]�$q��dE��=V���۾h8,wm�_'-��C�B}��s�nm�y9�2x;��{�ddn-�{��i@�A���o��F�GE��uR��QV��:RDb4��eu��Ir���i���������'u�tVd#"�G:3�
�D"�gʦv�~<�}��t��a�-��]C�`�su4��}����#>��,��r�D��
�"�R�]� <f���'Lc����g���iMY�HD\WzQ�x�\IN�If��BLk��t��ɟM/���Nэ�a��Td�8�ѩnD��>z�'��'��x�8T�����Գ�ɾ��F�
e	i�Əo�.�~���E!:��Fa��0�n�ȶ=dnuD�Qܳ]<����
���i�,^& ^��n#ܢ/�Q��:��6���QU�^f"n`hG�*�����]?P ?S'�GuA�`���i,X��z�%��'��A���^e�,�����-�N�Շ%v�f۫h�[x���`T2y�G�hU����!��較�
Z�H��y������Tq>���k=���V�JXt˦���}��t��ќc���瓬vR�X�ً/���]L�('�wO�*��3�F[y���*�e��Xc�}ce�E�D��ؐ�
��O6ͩ�~��p������SJ�h:���� ;:�6�_��~:�:/(?0�CU�j��y7��"�h�?A��5��F�b<Zd,�2BF0�7�ck�
��/*�)�:�ݫ�lg�.��G�PCp	lҲ7z�&�rv�`0��Ӏ��-cA�̸^4JZ�1(��<�0�U���������s�e^bAў���A�����!� x�4�v/�e�cW��:+?p
�*�7����?|�p�Է,������V6��,,�����Ux�s�/�v�ʬs��8�Q���%��̈F��X'`�旘��t�}�����f�<T+�H��ˏ������w1s�{���.@[:��Y�BM���Iڕ��Ĉ�����[袒�!$�?�!^�.��K�%���݊�䣚剔C�O ��M*Z�"��x�ԩ�x��4�WTy"��!��@�w!�s���&x�CW����_�iE�q�D.�I���(HD>W��P�k�\6% )k��뮌��Sػ���ԞB��8{�:����7�9c�P[~�����C�Z��H۟�~^�.�][O�R���=D��6I9�l��$���wD�N��9 1$R���LE陔���K�t�����&PI�V)���携{
g�	B�����Nj�f��f�i��j�Vy������¬! !e֦&�V,��L��UV lKJ>
7'l�(�j��o�3�~%�s_ �� �.�BX���cu�:H��ytG-�߳���e�!\eV��L5XN�um\�E�|5(�1��ԫ/THj�� Np�*>��;,��MF:�� ��5x�>������UW�\'�M ���7�Q��
�!�K�� ��`iT�<�F2y(�����5Þ�b�	ly֞���_�����g��7�0��I���G�A�0	@9q/�����0�W(C;­�o$a@�4�*h/2��$e��KdY,1&��O�!�D����ߕ#�'����AGH�Y��q���N���:�yz fl�>��z,�0���$:4�f_#O���?��ZT�Q2�xGl�-�E��1ʖIB�uUjNz���"ь��s���E.*���|������9�7�P0�ūp ��~(��tV@,�>0:�ۗ�CM6�5�^�g�7X<��X	���R�ݐu4��;^��4iDT>I �`"��(eq=���o�%}.�g7Y�o??h�b�����Xȵp���9o"K,�����e[u
���|��R&�������~ɼ������:z�D^��
H��hc��~|�[���bQߔ�6Ő�{��N�wF�Z�s��Y�z�R�-N��'D��ށq�SLrH����nȊc���V��G��3V���~o'��+���|��#��(�������V��	3)�-C��T���RH��^M`^�.������0�r7Z��ؓ�d�';u:�堔��1�y�C�!�k8A�\�N��_V�P���w�������� 8N��HF� ��IOzr@�Y��42P���R}6q'Y��
���3��Rʏc���e,I�c�0޼1_�Թ>������3#%[�e��?wj� ���j�<+P+w���|c��x�	���'
"�U��*r�~�o����	>OeOO��b���u
p��!2����}9�#���6�ALC�����z܃� T��I��WYaN��)x8���샑a-�����lv�譿{-�9p��6eK!m�����`n{�6kch"Tf8&I�,�qX-�X����f�lV���j�#CC^�+����Nrlf�;+���`��C�p_�DY�w�'vſ�W�ɹJu�$�P�9�pBɱr�	�y:x5�H��Ho�_P@�__��5CU��(�������2wBT_����R����EQ�ʶ��V�2�_c�5���G�\�|P�53�u@�۠(�Y�ܲٚ�>���]�]�v;�;�.Xi��ë��h���4�`f����T�.�*�<}:ST��<gz����֫��1�h���z%�Lل���S���P�����U\�
#3�n]�K?�T���\U$Fz<����Od
�N\���?�1���$؎
B�w2�j~�������q�ۣk����k�M��:iVG��_BN�AWl��
 �����{�0ݏZ��(L![;��Ne֍h��w1�J��@l��%c(q��^���(�
��n��+���Ddq+�hC�����iJ*Ή�\.�ap�g��#1o�X��*7��ƒ.|�x>9��k譳�g��Z|�0�RW~h� �Y�#��u�Z��k��8�9�t � � ��ll�}`\����c����7��Ak�^}�c��WEU��Q0�c�P֮���a9��e+:\u�J�K��%�;��l�KRzM�"6� GQ� H}鸰�W�F�a3����W��Sv�ut>��N��&�,W��{��Ǫ�09��} ��&C���|S"�:���a�kEc_姣�Q��&��8k��.���>C����n ������7yI��LM�뽢u��<��Pa����}�}Q�^S�e�|�$_���E�7g����;Ն�
Nu�K��8(c��1��1Rji�wP��kB��ǬTڸ�I�ͨ�����|�Te����N�6�&.4�.����@߾J�INԢ
j���Q<��%p}R&M� ������Y�8��=$�لN�@e�5�n�"Fgf_^� #�щ���A��RaMqf��/7��g�[f�_�Qaߘ���16!�л�9`>�D����Y�f٥�a�P��k�tb���/� ��QM�3�z�O��L1+�zh��
����On8 �J�Ct�R������:OT.���3P�f����GK�@�<��ᨂ������H\$b,ô�m��.����D$� ���6�@�p0��/��v�������Mm��6�.`�e��=i*}��p���\�M�l]��H ��3�$��E$NT� �/�����72��ɑ�R�y�1`�q��u=J�ti�`�X�V�����i^���ݎ��
�`G��K���	�~Kde.)��)���l���_�y�I
��{���YT�3�"��n��4Y��`�_bA�R9Yx�Bf�q�xɗ�O���� u�6�aƵ:39r����(�;���F����]��Ap���' B�P���'�jLܝ����",�[��7�x�B���Z����N�ѧ�5"��� s{��s��E��R�ɧ-�����,۪����]p���G���S�y��%r��O4aq�"h@%rnǨ	�`��?����a]��\�G:� �QөaĐ��F$��U�`�n���$�*���z�ȅ�f���9���}��=UJ��o$u�V���߉��z�����x��ޔ��e�����4���m-pw_*���E�SZ��r�� }WWw��K���%i���H'ߍ��G�����:�|yVsd����ӖO�f_��u�{jܕ%��Kέ�E:��{K��S[���!lK	s��n�ȵ�C�R[���oϧ�ȃ�y'�U{�h/M}QF?�"+:d�Ǧ,Z!n��CV���6yj;T黗�iҜ��J$�y��B�~{���2QZ� W[rp�rL�jY�t�^t)�|�T�*�Q�zs*7�y��e���#����vp*y�n�g��D�m3O5������3W��^�T ��qɼ1�� G������Y�U��ah���i�y�1�b\���h֤��*;�@{BB'{��i���v��5��5��'�_>�������������%�"3���k�ʱ����ׅ��?\������0.ךJ\���/*w`�L	����9��)��J<�XK?��җ�m����E�&�7h�x���Q����Ȍ%�Ϛ9^-�,j���o�����7������ƌ�L 6�Y�N^�O��0K��cB�:_��3d��F�u��0{�?V�Jf��+��%!�P_�?�{<2q��/[����kѲ�����S���8�7�O )�G��V��b��i�H�s��.�7("�.�/���)�`��hSF��ܢhM�[�~qo�~K�jX���B��N�+�N��C�h#��%r��2((q%ӝ_�M�lu-zB~Ѻ �x!~E~}$���TOD���g
y�q>�d���R�^�)� d��H�s��{}bJP��J����]�Q�@�d�q1a/P'B��&�X��U�`�`C/Es��?0C�E$�}`�n5����C�[����^�?��C�'-��'�7�ϣq��gv���3u@��f�dv��l��=��'��T�|��|�(���3�,;��1����1��&��_�j��kb�2)��n���h�	�$e�iI�T	�R67 ��e�ӹQ��ԯ�Hg;�m!��c:@���FV�h�u����u�6��]��o� �8h��)%���[b|m*`OM���ƴ�`v�$ɇ�P�F���A�98"�t�V4���y�U*)��2g;)ɽ-�e�@�5o"��Z]*���:7D�!X��a�5�Γ�o-��8�W�a^@�.�)v������ �a�ɩ�u=0P�:^�f���,�g5�,�XɞYMl3��i0��*�ժ���T��"������3���h�N��i�Ҍ/����*���B�S�#���h�ߤ���)2S0�/���C��,��=����i�7��5 �o��J�ů��0{P��n��	 T�w��!��a��Q�$�����
�z
��A8`�j�-����ḏ �t�v�䷝|~ Z�M��M������\�a��R �V���i�J9@��	�Nɣ��k���+ہ����9`�w����@�.+1R͝�E7��P4�-׸L.N/����"��`���(c���xe�\=���I-˟Ts(�)&�rId�H�|U����&m,ٕ�ƾq(�%��8�� =�ߕ�k!�4���'��7���z<ʎk?vSo���mM� L(�>�I4�����v�`��xkH��]�'�B�iW��*5!��5��}j,�\7�z���-�^<�.-�A�n.tv8���$sVq�C0�u�
}��C��ҕ�)]����=u�?0��B&ͺ�{mb���$��r�8d*�	�Fg��4���!*�a|&�k(�\S�6��XD�e�+��y�xp*��<r�����Ρ��(/�Ye0z40�^O<9����/���(s��=L��7�[ֻ�!�WE�փ��:A�g�L� �q�1J�����=Ece�Q~z� 0-F�Ǚ����?��&��F� r�����y�Ǆ����K;\;��[䈙'r�q�NsFd��"6:|{���f���*.����+��A��K���R"�#[^k	*/�Ҹ0�>�B��e	q�(���H��7�U��Ȏ�� 0������|&~o|��6����pWm����[�G&ܥ��[}�x ��I��@A�U׶�o��bX�[������v�v�ݨm�ݜ\HnH�����Ѥ�LS#�ۇ0��M�똄���{����r/=H��װ?ѱ��12Rl9n�+`ꟼ&֔�YCB�Ct�r?�rŒ��,u���Ry�Л�$�TTc�AB:=��|��~��r&x�����ߧ2�7Q�fZ�����x3
@>c�1����ï����?l�6�O�Y��0ئx�?ɩF����[.�r���k^�x;�t'�C������Վ��A��O���J���gk��b} ��G��� sI?�K-�;őҥNq���KiQU �w.��u��cleE��^-�w�E1�L��7�)�n�T��;�KRZ)��*���f� G�!8���ggog�n]���d�&Ao�@�i�'&�a�"��Yb� =3��Wb���M�*4���z�ˎz�l��,�i�+��Pb1�s��i�_ďQj�~�m:[e-������&%�:qY� 5�8GY8�GCu��Á���O�'���y~o	3k��CK-��c�^���$�m���T3N�%}��>:'G�R�',�ٗu�1��,�O!���۴�uNV��s��ޕb��,��a�й8�+ަ�!~U��0���L3Y4�CN�|_�|�㈔ț*�]iz�$
�@�3x���ً c�.��g8��]��_�G�n>�'@$l�p\�4�Ub/2 ��i=������vG�Mr�^��*�2��D�5E��~�ߞ<)�Q9�d�ek�WmB�hnjʱ'��ʇ��S�=���Z�I-G�uh���+SV�deu��F|��Ob÷G;Cn-����S��N~C�3];�;�g�+:�O+��8�=�����V�(&Þ\v���t�I`�nSm��[U3�c���7[V�Y1���Od��N%"b"]f�y`֕b����:�����ч�C�6ӈ�9�x�V0� � �ɪ����コ�*�&��y�2�(PGq2����\�ωD�������NP�Q��C�^�08�|�U鏮�iX���!¤}W|�
V�?R�TqR�2)f�﬒�����/�y:�t��(-U���؁K\�Hܳx^�rR�tS��r0y���SͯC5Ɲ��F�/:Sy�`��B���g0C�8��R"H��_z��1<2�ɷ.�f�@�Mj�]��a��-hS<G5f�yG�? 	�r��⦔�;�E�K��iT����t��A���=Z��G�&e<�}2�#���N��?/N����KBp
����@8D�u n�j�dJJD�;�M�w0A䞘"���YF� NrT|Q_|[���:i�H7�էˏ��'nF͹�������q���x9ݮ�(,��h�3�F�ۯ��I�72�Fњj���߿�uAX����]]�<@5��o��E��ji��hԇ�i��i��e`��_�rgB�����aO����G�E$N�EA�v�Q����a��Ӻ��Ʀ��j�s����s�S,�G�t�*����l��>p�@���qv ��<@��~͈�	|7���^v�I�*�{�g�w�fP���0��p�J�sE����ߔZ�9�-�A�p�B'Q��x���x4І7������.H�F�9����u���^Bn.�IY�,=,�/�{����ĀA�G�C|�rB����X���Jd�,�}S���PSd[�1$|������P.P�`&"j'��#�b�m4����W�m&��x���~<n�樍���l(j��BL�]��
,�
W;����7�����8^����4.0����������!V)�6��x�U��B(���Y�G�۬�͊�u(i�s[ꂧ�8	DX����4��4�S��64&G��A���w�k�����t�xu��9��$"No�'�R�+�NjT�7��1	��9�5���m>)�,^#�r�yj�#���n.�����n`�7��Y�o���
��(��*��m.,��J�D`z�����.�{�T��$���践m��6�Y��ǰ�beZ�?^=��A��̻-g��vJӐZ�������0���0�����)ނ�r{!��׊_��3��J&\�I�h><�����W�6�\X|y���[�3�)~��I4{]�Xg��"W��{�PZOѼ�����-����y��ͧ�y�/�!}�"<�n�V�P8�]~�A�[�A\��ſ!P�@W��$��K��:Xl�]?G�B�F:j��Ds�B}.��H��G{8�;�����+������߅�DӼfh��D�lm���������+�7W8�.y{���R�b���\��X���z�_~r�.%��~x�ö��3-J�.>K
7�@��1�%��E��o�}֔Wc�OE�4���qzY%I���M�-��Ҫ�fm *1�
~�*2\�Zʡv�`!|s�;�H�q횉IuߐDQh��s�mk(S �{'{�&���а�� �҃�y|�X�b����Tz֙0���5��f�w�zL�� �a~���ů��TDh�L��4,Wh<���E�"ob,���[����i���֯I�6�#\��8{ӱ��&�#"�#���SZ�C���	"��=v�YQOC��%j�uA�	�E�wڋKN&@�~|.jG%	�\'��E�X���[�uF$9PH.��a�ds+���_G�
�~��Z?]��yV��޼r�O�r�-�G��.!�����$W>M�_8��Nυ&E.�@�S~�D\�[�e��>��$��y����o-�hI��Y�q�8�v�ݱ��uw|H9`��8]�S��Kj��'����}G���3��]_�&��3;χ<����K��ŭf���@7bbL�dp��е�k��M�n
�3P�˲�*N%��8�i�l@�z��U=�]����1f�,t��|Ќ���%��y��V!�6�M���W�͸�B	�"�~ht7ݩ���r�J5ɦ�0�~�:�A���e��`�t�����@�=�"�Yu����T�2�[��x�|�HT=Ob��B(�x(5ү�g��[4�5��w	�.�&�xw�����T2ױ�W��wZ�����))�����{�5Y�9 �1�o�1А;`����)iO[�+��,}�mT.A���-:9�|��b�Vj&��x�ߔ�|�B�ȍ�Ĝ�4���"A�g�m�I�8+Ƽ��p�(9�1m#?n8ɼ �Ar�Ճ.�3y퓨k���Ӯ�T'yi�s�(�U�d����u٭ђ�*Bn����u�����[�\�.����ˈe�G���`N|��Xr�������ԫQzbC]�U��-�
x 6,� ��7Ve��G��7%j��0BvƃC&(�[�]�X��.R�su�.�B�4��g����iE��S!4Df�������؆��9�3cX�Zh���TTbm�䄢�Fҷ��[���JE_ģ1@$�o��Z���������[Nn�JV�T��I��ㄊ����Iѭ��N#�9� (���>��d��fl�r��E񶕴|�UB�2XG�!r�z^�yU�x�B����tf��9W�K]M�S��3B��NybM96��K1#p���9㘶g�Y��c�3�DG�-k)`�Ì>�m�V���
�_�L�k��0[b䖒��%
XP�$�E&l}�ʬe��Y�/)� �9cא��˼�-؜��m?������A�Kc��b��U,�|3[��C[�N-��v�Ea�A�pAܭ���.-����3"&�~3@a:���4��+vE�y(c�t&��e�2��F��r���ՙ2Qڍ�S�k�# iG� ҷ�=L���:�7��j��t��
JA���?�c��	�/��D�����#���+���I�B�D7VY��3�ז�[J$����dK괘�9�(Q I�{��l��S��cI���]��S��q�����X��^�ǒ�6^�\Af����ui���o��m�f�	����E��,��a�ޯ��l�u�����)�	�JjtW�2�%sC��v|�I����������ozC�d�%ր�oD����?����>��|�	�[W��Z|�!�����e��t\�!��c|٢�L.��F�{�4p����]�.z�g� 7=��Q�=q�^�����Fx�����!҇��v�S��<���� ���n�ԁ��d ����r�!E[J���r�Uk��kE͂ �RȆ�K��J�d�{eUx2D���f�T
@���xg��:=�^Wpndsn�?�f!������X��y�W+́��G!Q�s���qM�O�T�D�#-j�BiL����@g72�<D�R˺�X�9ފ�[����\@>-��'5�b�Ɩ��ð����Y�e�X/�FQ� ?Q�K��%I�K/��Z�e4��9��
�����U�>����u�  �&4�v]�t�H��NV����-`-u����T�,&k���,���b3o4�ʒ~*�w9�W��d�(��9�,�:�o}�@��;�0�����O��-�T��2`��w?a��sVȀ �B��w� �v��'O���)�q� @\-���TW��$n�&B�?�+{�5>lP%�	:�%oIM�Ɲaw>en�o���&}K�&-�#��q��ma�Ą�y��Q'B���+?z5y�Z۞}B���0|�GS႔�t[���Jp`pN�.R�`y1�㘞Og����F�P�1(5��&�N���i���_C�P6Z�wٛ�
��f&��En�!��ғ�1f�8H�����8D��W5�H��AE�QeP.�k�0&'�5u�K��*�ڽw�@�;m�Qde9�(��b'�Y�O���H=��F����F�O��{$T�W??.ցa�b�'�Q�7ת�k$2�'{�i��pJs	L��x����"1ǁqy!;�����@�$6��!_�Y'�W�.�pKfۄ��xU�T~Ү��9��n����2)�2��=�^�<��S
FQZp��%8VFK[��}Ir�S{�ʕj��J�h]0��M���,嘏z���֍F�d*6�dIh����wu# <�Y= ���<ᄀc�C	~MA[q6T�l�ӿLp{�ٯv�*"$Nw��luǳL�fR����~-���'�X���	{FyyK�R�gƸ0wɖ\�^�"�[ݴLU�Atn��J��^.�DNxa���j��|��ߩI"��`�rI�7�?s�OC~��e�I�]�|��wa��k�m����J��;h�hQ$�V+��({���Q��X��R����?����@ӫ����CѲ���c�(��PN�9:�|�JM��T���>^��	c,��h��
��օL2�0��f��Nu��y�ޑX?}�c�9 ���L�ĨpL�=�AQ����a�~-0ٶJ�4HqDOv=�8K���^�3��ԤB��>i � ��4��O�����Z��Y\+E@��� 7lF�7c�Zv3�����)�S���C��ДC�^	����bs�HG~����������,�S|L]E9����ҩyUE�=��/�Yf%)����dm��	�	ٍ�"�!�ک���/�c����̔(���ʡ*{�O~�
ϟ��* �>�"�i�tI��xȋ��2>늛9$�Y>�R �ŉS�?r���p�1K��^�H��۴#��1)���
R(`0�Wﾶ�ÀT�$+�}
��9�H!D�-WG�e�S����F���v�I��PIG�qT9��yg�I��C�"xQ�T��ɯ#[2�k����g�GQ<��T#Cw�;"ņU(�e3^������v{�������N�bH�n��t�|ݘ�{�m8��T6�^�t�ɬ
�I��Cf�����yS��Ç�ɦ)�7BO�cE�U���]��m��ӵ�/���B��,� ��z��0����ytu?cĿ�c�x�NQȩ�"��x0;t��S��L##�V�{��������������6�5J��]̀�bo���?�������h��"t㙹�BVDD@������4vf(7�&��h�O�����z��|XV���5�a�����.�y�#��P���� ]~���a?���}�ݾ�9L���e��d���|�:��ϗ�>��)��i+��;j�PĆ6��?�����kWO�?��~�cS3+s�W�P��[t��я�YR�x ��A��Q.B�f�0���yxZM�B�L�������Y!��:ޞ���P3����t3&�k�ر�tށ�7"�w��Ю�>���9SSI�3W(w�LJ�mIp^\=��ȟ�_�������W�m����MRy&�Y%r�5�D�v�7��q���.w�|>^ږ�^P�RT�a�j�z`�^H�7_I��ct�š����nep-cn�@Gj��BUM��[����Zk�7�����R!G�;�ը-h\�"{�҂��W�Lg�t�N��NE2`�T󍫂�ԫwS��N�A���ZN�m�E��ŵS��/�I����+Hqخ���0�x=�bJ�_YD�E�W���!�z�t�7�\��|縗�@	�Ņbr$K!�V�$�QR<����>�!���z�F�V�5�jy�|���j�wf��P�D3v�����g	@��-����&(�,�P���OC�q�d�Jsŗ~�S���c[P�b~�Fa��eS#���CW,��S��^'�m�n(�����6qZ�17�t����bd<}Z*���q����6����>ژ2K��W���^Y��j[�)捊�D�`��k�6�Yb�l"���Mኋ3���P+���y3�ʛ��k����P�1D(!~9�a*�԰V�>:�OaY7��h*�6�Y6D4�$�+�!�S��u����O絇�\�NȻ�:�x��3W�1V5ˠ1���/F�63��=�,Vt�R�=E}8���~$��������eKBs��L�1=o�&��C����>=u�If�Ώ�vip��0VXXQ�A3��ޏ ��\eSMC�{l�%���k9P�FtA뢭���u�7��E2~�Q�U�Z��w>���QX"j�`�A�h؟�7\��6���r�)�"{p����c��)���p�;�U�A��Q��@i��h�l�_V�djR�YHX�PG��t钕�d����ᒇ�2���M�4Pd��X�Wn]���t'O����i�Gi�2\��nRzsG��?l�Y�Y�f�X�{�ӼR�H�+=�WƍT#�mEIYǪ��$��U�M��~"�1�$DF��(i�=|^ 'Q0JW�]�W�ɧz"+�"N����j�WP�}����W�H�D�\>8���z��]�dEfI��ǪaM#�c<A�-�HB��W{	}v�RT��Aѵb��[�	�(H����n�h[���"+�E��XT~�M�o���^I��?a��I/�<�������"\ر����V�pqbU-�3��S�{�DW���d��X̚��E��(#�Ns�d��4J�G��t���'GP�
MF"��R�yA�xh��#"���B�Z)
O��.�.UFR5.)���p�>�QV�),[8�|֯�uJ	��Ҹ�Zך�j�(v�g�Ђj���A��
�>*��D�j�G3.���{K�ӎ�@@�z��"��R�1rk�;ķ���YUQ�7��{`M��$�Y��n2ű���z$<&p�rV�K]m�{ְ)|���SN-D�.��]�~K�I��H�~ה�"]"`��,U~>�L��>�)���/��Եg�K'�a�F;)�k�=�����Z����l��X�T��x�G҆l�2�Ky>@�)��A�����rS{%��^�-nW���gY@��x�"l���hq�pĈ��&Ύ�p}�r�(�^$�o0A4
	�C۱�*��u)��n��Sܰ�LKhVEsk"�&�"���ݤ�} �X�=� s�Z5ͱ*�V����'��eJ�F=z᥂��)�Nҙ��+)]�,�E��<+/j}�=`�ؑw����.��;� i�4:�2'����J.���B�k ~�3KB)8��~�Fŀ�fz��.�h>Q�5�dI3(�X������D]�	|�~ٳn�+sO��"��A'�%@���&,�n��Z��o�>O/�P'�b���.�����H9�p�7�k���0ٳ���<�|�4����Y�����+�R_��>��fAg�ozU���j�W��P_��4
���/`����s�(+��9���:ԕp��S4���B���©x�$Lg�!��h���+�8%�ߐ+w�G���;�i�)�	l�g�8h��b؁AG�9�-z�ߎe�qjl�0��3�Ԥy�>-)�\siH7��p�n2�y�0���!�&�d|Y����Z�Vħu �����~+=^�u&��:�޽�aF�/畆�2���?��-�5��M1@�1:��Y<8��E�wy*F��p���d�h�=e�YIA%�Lܖ�\[�������"� 0��k��)s�O�Y5��$��0��g$��E��_r�#�L�U�#�N������!Z*���>�T��jF��R*~�K��W�veCǼF��fqh�D
R��R��15�D
�pIx����V��T���5�xQ�rO��t�F_�=�f���"�+�?;F���o�Z�/�x;�k�k݋eJL�����<�����ȁ�)û>?�J�͍J飒L"D�"�����Ɗޫ=�^�둮p��D�hI�e$͐��k�^�C��4LpE��j&;4j�y�*Ef�iR�4����� aA���ՂXdf��2v!�Ny;������4���f����Ɉ����Hb俼����rt=(r���6Nec�U�l��2����,�JuA=�m��<eV�^��]=�$��;%�4Y�t�R��
���	�vV��ޅ�m��j�@�f̂\Gr�����\�j�L/���v�|���1� �w�F�Y�hX�	��j��Ŭg&Ź;>����ٹ��<*NO�b������	�Qߐw�,��a_J��ш�)W�tΞ�U3Pe��+3Ut0_�a�������� �5����TNl{��~�T3�4�b�X��P����&s�Ƣ{�W�� �f�k+��Z�|	/�e����b�LZ���bh���Ѹ���*�;�+an�_ё+ƃ��� 0̽��*�Q�N�����U|ϓ�^t+� XD���n�j���#(��ݬ�D)�R�e���?y<�Z�5X[�f�0�5}c��t�:��l�5�1v+YHV�8�.5�����*��?Az.�bmQ�H.0�KdQ?Ӽ��<]*���� �ѷ����ݷ6��72ap8�z��6��e�{Vrq��k��G�T5���P�p�T1[vFv�yy��4��ߏ�����'�t3��>�%6��=|J�w���B�j�M�=����N����M7��.�S �iP���ўDk���3*.%��OE�t9��5�]�h���x��̈́��Z�Ǎ�Vhc#�/��O��^L�Oo�D��~��3�3�=�E~�o�.�'�}`��V�6P�v��	�3U{>x�!��^?tqe��()u��J׋��p�0g�5�r'=æ.��`ӥ=�������_fŬV�<�%V��ě{�'o��Wz׊n�e�u���X���zF���KH��H85���)2{X��+���'����/� I��a��`b�:·.B�G�]0�G�R�!Pp�(�ɀf��e^?O��%M(�=[ȣT6�I�����<gä�-&�>�׬�_��bA��:S�N,)��	�ư��V�P~M.J63OH�-���-�C%;����X���g����q��Q��!�ӏQ%-��/.j��/�F,Q����&��ʂ'Π��s��P�;�|���,�%��
&J��@�R�ڨ���I���h-ީX�'a�2��d;�r�~κp���{q�8�ˤG���ݧIß���K�����I�e��J���!�������k��p����U3� dàP2mn~BI�M������騥>A�nH4��Ҷt��TdT,T�Q��zቸ�m+{8c����cF��������f/0�6�3�9�w��शg�a���)@�������P��{�� �߶M�'����!�P��,YܣU�|ځ~Muu���jq�rpD_M�//WK1Q�K��oXMj ���ǯ(�Td{�J��ً�B�
U�F-�`�z�Q�:���*7�>�Ib�Њ9bZ���ِ�r���B'�����o%��]b�ާE��tm.�����XL��EI�`Z�����Ŋl>Կ@�'oBcN��w���Ҿ�ĝ~�i����0��1਱��.����@��o��t�n������25ay{��]��Ɔ�1<b,�-��ӄ���共/Մ�82�-TqAD�|ÅL�	}M�i˥�ı��q)�PV7!1�o�xBY�D��ⰵK�̆!���|��G�-�8�\�'*9�O1NN#rX^!�
;�\{��9�&�� �,���uG�\0X��,!��>+���}���ْ@�q�L�Dmc�>�kx0�R*[�Ģ�w���Q_V'��Ӓ˅���N�EP7Wd�G@b���F�D�>�����2\���VI��U������:�}pc��9���hCe�N#!�I���o��N��#����CK�F&�		`;߆ኂ������LI@���:`��2�A��!6�U;ȃ�9:��_�=~U��Ȋ�S��~�Z��GPԶ/�L��!���ԟd�WQ�2,�|x����y�ݰŅ@<-�ڨ6|�CY��:��|��է�IpQ(i ���8�G'�l���,M���0��XG��&�V�Z2W�y[K؁��ҹ0B�A@����czgeh-l��a���``=��"V��0�ww-0�_�?��S/��Y��J�߫����Z�m���	ݎR����R�wm��Nn�������g͘�0IQ���f�#hN�L&0��4�z����x�`6��]z�+T����K�=yW'�'e�Dp+��d�C��� �d[m�h�,�gy��,�Rbթ�K6��E�R?l�n�kW�=M�b�:�k���'�Z��L�ъܒ���e���y9s�3�s2�$\�����'@��ZM����{'G�3r�Wd��ԑ�e��<�c�h#CK"/�m�kb�`���ݼOgB���_��Y��4��jQ2����{�c��Rԯ�Zt4q�E��2Ʃ���2�����X���[���?�v���E݃bˀ�1u��+ĸ�c�WB>x*�h���q�̤�G�&�g��RXjB���7v&t~&:jJ��!c}`
 ���h��� �_�J���\�	2�͆%Ô�[��YО��Z9#�]-� �!Q���N������A�G�i?-0�*��z�Ւ�"F�,5Fcf�?z_�=�T�c���'������ �R�d�E����0q�fk��2�Bv��<�o��^�g�Rh!�r_����0�#�߶�"��M\(U�Y��g���Tg(�C�k�ݥ������>�Rh���[1[����r
O~����<J��\^��5#��w�S��b	>��q�2�L�b�>2�R���|�p	�V�ߡjz��J�<���4���q���u߉�^خ��+X���� dNw}�G��_�AB�I_��o��_����~�!����!ʪu��Jt�����S��q�$L���5�؂�����fI��ţ�M�W�������@��ݺp؏������Bɟ���-I�
�A�O��+�������2z�T�g�P&"?*o�5�PƯ�����:"?��TF��t�'��������םS�(�zg�+�z�q���R�q+�k���c��t򚣢� �om	4*[e~���X������c.��M�b�qn`��DT7��&c}�0�����1vȄ�s��Y�$��M�J���,��o�֓A�ڎ4�Ma��\�z16)��#&���3�tU��U
Lՠb�pT����ۂ���B�CwL}�rY�N׽ҥ#Z8sC��&���k�����z��?����;��|&��"�?�:g��d�m�A؃K@�Dn�����5{�s�
��S,���ա�-z�[�E���Ϳ�������U�:6&cxc��J�kK�įr@t�Bf�YL�(��>W[�R�2�
��ߨ���K�ΔKܟn�����`^�����k�(]ml�Y
�r��!�?�H�!�mH`�U�
��|�!�)'ƹ��W���fXJ�����K�ʽ^��kq�J��`o���)+}��p�ǽ2�����ĿE�J���Kq����L"��\��������DR�%:1|i A.E=�3b��R�
U��w#9HV�AU( A���"b��3�T,�g3���	wu�v��j�ko.E�Κ���K	YT�����(�p̾���+�S�1F~��L!}{(��]iZ�w �AS)#�6�t�9~��*�ku��R1�r�%��@�+ޒO��_��r�q�n�	�w��i��k	�����M�]�v��S��&Rԩ�-C]����L*Cy� �(d�~yOG�M�`�K]���+.�h>6��a@��_���&}���.i_F��A��#���T�h�9��R@��~�S$e�����.�'E�V��f�u"։m�f����F�������_����ZJ�C3"-z8HY����b�� ��hM��*|]�\��w�Y�,�u0���a'q��ȃ"Ϧ�tH~�!�K�E}Mġb�._�9#�dp�X����%}4�(�Q���je �d���Ce��39����6�h-
.�'Wa���̮�{�+{��	��u(*K-G�#Z�(.�
N��8Q�x����},�(:c�A=zdu�/��E�@�
���S���FI�Ih$�������O�yA{���(Zh�ą^⠩�04g:���xI�b@��%:^m��sq������=�C��2��,zQ����4�?�Sr+�Z�u������fVk*��Xp�f䯲%H�Z�ѧ�j݌�֛ɠ�B����%��'��tI�\�IA��+^�fi>���K� A��ڶ�F�x���Z�|t���a���
Ń��k\��M W<2�"��D ����\�}�U� ��j\��@S�&z��\$�o֤ZPܜE��r�1��
�GS��/���Z�;D0A}W;'\YD8{e�h���R��C�h+Jy��+��؂�A�R�V/`�*y��\˾�j,���B��2y���V�ֺ���6%JAW�F"j'�����#���J���@�0�G�t�!�$*�CxO��}�)z�o��l��{dNM�[��EtH�q�	{�v�D���c9��s�� ec=���C��R�5�K'^�tW>��Q��CD�?ˋ�$Y'.�]t��?
(��TBk��B�,�~�L�F�Z �x�(�(��>2ӓ.7c�,��x�'��-tN$��8\�aC;,����n��t�e�h	Ûf�o�]]��.-��4V�2��i�2��貦�x����er��q+N�{<����9�|)�[y���]Y�Q��^�T���u�~W��:������G7dm
KA:o����O��U�f2���!��O�⛎]��9�+��h{Q��U���5�z�K�N��esԘ�Ͷ���D�h����^3bkэi.�����N[�)��%LSD���Ta���5F�o�DǱ��ٳ���Ҙ�C����pV[P�����p���e"�v�q=�Ϻ�V*��?���&�_�) P���X��K����ͭ����/B�8z�7fk�U�m�,�y���{�*\rŞ�P��� �P�|���fe�|���S�Q�!eOR>��}�N��K�7���r�\ /a����P�֢�v֕�D1�W���+���i�c]�	&�u�`�n����t��j��Uc2���j�˴+<	���A�#��k�1N}T��ڒ��ft���2��R[��H�����aB�H��϶$ď��b��E_�wa� �K��c�5��fZ�R� O�۽`=�	خ&K�	�'��6�ݑ]W9>�>Hd3\U�D�������gxq�nH蛫��醓�E#����7e%�C��3;3<t���kLc�<M5H0��w<G��?�32A��PvT��K^!�H��,a����Z���k�9?��U*7�X�Çxu�_�l�6x��u�8�Aմ��ڽ�K�:V*=F�U��	��ă[[;M���(=�X ޿���P�3�5����V+Pc���ֽ���Ջ=�ƅ8.���\s��@}�6fBI��4j�+����,��p����p�6��`x�C6�^����(�q_�/?Ə_w�p��Է�4Z�<TH���/g��G����2�Q�f
�Serf��L����S�F�rJK����)�׊�Dxa�����)�*�oVX1�����\
t*���(����n//� �["����Ad|B��sJC�$���U%{���PnZJ�X����d�Jk�D+-(έ��z���<#�V���. #W��^�6pB�=��Bw�L~��m���unm��1ݕ��#+O�ˡj���6���wG� 0!��!oZ����[w�؀1NAh�*X��P��+&�گ���c�=�[�����G��8� `�I�#˹�j.�����-~%zw�R���U�a�|�e�Qw�p���D�J=s���89��G5��$9��y�;.}6��|o��F�3~�z�X=�9�kkgȎ������s��b�U�\��s�^�4;�Ӑ�0����)>�_M�Ga�J �Z!�W��m�zX5U+_a�\��8߬�~�ryH� �:����-��� S?u�PP�I��	����=��$f���a��BQ��[;T��f���	�Nce��������;M���4)%٧n�m �nʍ�,���0�p��R��R�NWǾ���؃Ep6DS��/���HW�O��|�O�wMS[h2�Թ��C�51?�%��@Ɔ#%�f����h�,��}*���w��i�����o�q�%�q��c�e�V���m�*�����M���Ѹ�p@#��"����t��&tmDi�t� 4��[������*h*C�#\�Sjy�S�����Po�`�Ӹ ��O��*(��]�P�v�Y�U���$��H���}Y����:���/a�N#}�>���'��!~bc�	#�e@Ss�fܯڬ�yv��{����dh�l��E��6�c�>�G��a�M Gӻ=8���Z���GwU7�p�-ϻ�E�Hn�����fS�V��7��f�x�᳔P������D��?Z���rm�F -8��@��=DjB�m�TzI<揿8;^��> z��ӣ7&x��ȁcY��X2c�)̽�_Լ��FX���ikT�z�^��L<��L�C"u偡�څ'�*�iEV�e�SkQ��!�%��[�œ(?�|6 5oO������]̜R�c��z�z�F��a�-csZV��_.��fAܮ.".��I�hk�`é7_߽Q�Q@��ȺT�;�c�*H�+juOD�^��[�Oێ̡g��?���H��}��@�z�GlҢj��-|���+L��W��2�(�xl2��vAx[���r�2V�	a��f��=	������}S{&���w�'.N9+�!Ҿ�%#�*�WSG���t ���㕮"�)K�h;��tc9��)�M0Xv �w5�즐G�GCBI��4�A��5���p��м�6��ȅ���JΔrK"n���66�c��k���ӳf��#��F�:�1�`|M��rbe���g��5�Z>fxX�c[�a�_q��.k��I�bE���0���r��VIb�ス!�>��K�qqs�+-�x/�
�ey�g穽��Z�=��/$�|��f$���^Y"m~街Ͻ�|�5tTCFUq��k$�.���b5i���cM-���/o�-F�\s�+k� �f
��	O0��`��	�Se��@*�>Ϊ��_ֽ,ń  z�Anm�آ��~߹�5v�����'�&_8���"J&��M�I��� �Z��_�x��\W�b��\\���l/}���
V�^����G��}���Rk�������$�1V�έ"�]1�!������R�Ʋ��K|�f �����"�е�|i'1|F�6����Tm��YE&�1�����D�� �H�K-���G�M�z��$��"��WR�eZ.޿ԡ-B�*|�������AO�m��tud)��}�5�I�pQX�?7�����!9�!�4��ߥ�&5B1����%���c�}MΜ��w��E˳��<7,_�8M:-5k&�/�� �/O~h¿���{���Y����f0��c�'V3�����F�q�F��=暳�����V�HL)� I�i��zE���r�WM�,z���2��4�7P|L�gM�E��#!���ZQ�]@[�X�U��޾5~��FE�P�4�~�g��]B�d�RT7pr �ܯ��X��V�7^W�����N_��VK3�b�d�>�<@f����c�e�٬��kݛ��n���L�B�WEI����ݗ��"^��s�M�m^E��,#6��[VN�f�c�@�*�Z�2�$]]�Eg��S �V��0����tr6�b몫��K��]����䐪#����	X腷rQ�H�OǊt�Cn����~3�y.�"�Kˇ.(��m�{�fU��P�s?}s	����q�W�Ri�Ec�<�D�TR�@��D�BP�����x�����<(#?��l����9��yD׸�	Y�ߕ�kl�
�ʓ�q��t�a�1��O�=��-���RHW�ְ��,����<5:W&{3�&���@#""���##Bi$�F2�4�:(�;��Z(��&)p��<QOI�� �&t���
3l�Qe/��a���,��L�e�V掻����D�rl%p�t�!IT�G�oc���7�sU<P~�Q�w�����dFԙF�p�/	9���7$/�^��>��j��L}Q�qq����l�<�<�yI��:cc��62����S��1�ddD�^{�B���?!C�py�@Q{y
�����Y�kی�ӉZCk�<���70��|!>�:x���\��m�ӽ��v�v/�ݱ�m��J�ğR�Ȝ������(9���K^�3K
�9\��e�ƺ�7�{�K�/t�����;�QL:�S٨��nɔ&�Y��"�P�W'.����NJV����,�p7SN]��ҏ$��F��E����b P�>�R�<���-�J�`&�b =�q�������o�J]���5]�բ��=��@�~�3��1}?���c^�YM.��9� e��wο?��i���p(���{Z`F2�j�1pR�'���	��*!s{���-�٫!n>�#"��aF�����Ό6ɂ�9�@�PO��-�66�n�����3V��ګ0�2�A��֡��uk�Py{;��֎!��@�eGXV Kɭ��������7��e�#�+|�I����H7��ժ������_��x����"yW�B@��_��d���k<�K�����54[��-��v�L�)!��Pۧ�v����2�wH���a_��>l�B+���A�R9�:�W������� Ta2��:�>��������'�kZ���+D�bq�I��˯ey0ܓ�C��Tyr)�C�;�W�a��,��č^�W�Ə���p|}�熰��������t��r�'O��s����yHP�U.p��.L�j�slʎ����B4G���eSo0! tj��3p��(��4v�Ϧ�b�f3Ah�����2Rg��^���\�$)�F�#!�e�q1Z�?����ŵ��^<�̸�C(��j|�E]H��*W�,���s$Ď�X<*�,{��=oc����P��V�ܟ�t'����c|?�&03�!@h_�55�y���C)�᷄"\����B�]�X��c٪Hu\V������D��{\�#��Zښs�CU�u��G�=q�kλLN4����i�@����k@]`��,@���E �.)^�O��n�����$%l��L���!4� i8vJA���]_�֋�q��<��L�bw,��o9� ��(`�����'�f��~��@ �����*f�θ��7b��r8�q�0J{5���.����F��,{Q®��S�J��?�qE��� �\�F��!9�QE�I�*�ʧ�Z�ޒ��U������3�"�6����F�RKB�3�S#�U)#Nb�����O`��Y����e��
���.5Ɣ���A��D߈�x�!���#�^0���<D�ċ�}�̗^&� �:5�\n!���El_���F���]@��x�:+.�S��fb��E_[�S�q�z&g����k������U1�����D^�R���fwKT3|9`yEȍ���~�n��<;J<^�ػ�H�]K�C�-y]p��@��0�n��W�6�T9�G�%ꝧ׋�t��*`������!���]�Ᏸ��c�_�F���ffn����7s�jf���1ai�X�����dZ&���I8�(Y4�T�&q���"�$1��a������qd%�ϟ�]�j�<H��Hi�ݜ�.�0 }�b�*�1u�q�!E�d����؇���hy��'��^�̈z� w����~�<��Jw\D��\^�8��_�:��z�ξ/(8�fy����/�E)\2���<�}łX�^�3��nlӷ�B^��u�`�F�BI��ﺡ�u��p	Zh�)�[!�%�aE���Y�=�17P��m!��̝Za�W�E�bL	���-t$�I��'��À��/h��D�`��C���qW[�]U&��}۰��z�Q:�����R�%;��ϳ�~�)�qG��!�{ܱa� 7E"����z� ���.N�/�����ɣO�<P&�k�u����2��$*�lw�"1�#�n��%�Ԟ�$�unH2���6��PdQB%ҳ�ֲ~ާ4�K�,�j5��kgх�X�:WQ����.5���d�[·����H7�����!��Ħ��s2��u��
�"�&t!9Y���L�/��S��X2�$	}�����|
��> o�T�x�������&��	r/�#�	1��z�%���lB�{	V�s��'n����(�ÞXG�碍A��5LV�W�*�3�t8�$�⢔�eR���������n�0���[i�M���+iĞ��0b�p���X$�@��_6���	��[C�ǳ��>�O���nL���-�4�\��d���?So��m+'��B�b�y��F�h����f�Xۊ�����o�s�D悺M-6�V����|���q��ܖ���ݝX�eR	�����s?\�3;��A�T�X$�e}��e��n�ž�U��PzV�_���o	;_ұƼ���}�f�j��H�
�W	vE�À5/��i ?�$��`�u+���ۻ�q�s���1[����������Z�G`����F��G��oy,Q/jbĶ���@7����K
��4��"�K����N"�,r}.t{�3~Ď}�Cy��;=�<6͟�#O-C�
�qȵ���j	~d�v��0P8�1�,�h�n���b��`D:@L���ۥ6��,@	�ɾ�}�1��#���jV��[ ��a������{�pcE�3��~PC�R�ɒ.QI+��o�s�����x�V<��(�-�-g��.:(����]���.��C�0�ݿ�Z�]6RdA�2&��C��Ƈ3���W�u�]�G%nm5��mTG�gY	�y����ޤ��}��MO��-�����i`��ƙ����rxr��ᆚO��R��/ Un�ks0k\�B{��Ο�H�'ýj�3LR2����#�,]�$;a�=%K����`٧5U'i�4ZC��־o,e��Ґ�0�����@��z��w6�k���wKi�fN+mWI}�LX�L&�т1b�	YB\<B)��m��?�']Ís����vr�n�W�Dz�4j�zgnj��G$ՙ#�E�s$�J�{����|r�	�I&�U4'�0�c�9z%}I�P%�1p�s=$n�F�~>��<y����;�?po�̯-C��|�N�[I_a��W{X��B��|o����ąaoJGn^@�|�E0l�w�|�Y��z��U�}���1�V
�sw����'��GNҹ7�ۃ�}��,���\���W�z�!b����7��Fƿ�x��#IͺX��}NK�M+:(Z�k����Ô��9�M|�����6k�n4�V��+��sK�j�Խ��`�?��S��y�����<p�u��pPOUP����/С��S�Yg��W�~PB&��8͓�DS��c�LT3��y�f�����_���g�\���5�����TgY����c� A>�[f��g�,NYw��g-�[���?g\,�^��YSթ��_�
 ���F3�ﯹ@�E�/����w@6����t4D;�_���c��d}��^��{8���B�f�{;��E/,73cdI-Gv4��'��W�g��H��/>��,h�.�q�
�lƖ�j��;�0&�c�M��qд�J*�^K��~4��	�S����~�0{�0_�v|�W �AM��}(0.P�Aj�B�ؒt���b��ઔmx�a?�N}��"�M�#P0zJ��=~)��{�M�_	$������>M�
���Ռ8Rs��	a���ʼ��:s�v��%������������f��<b��S�{�P4�!�*�K� xt�6F���N/Vp�-���f��r�x�Y$�2s�[FE��4r�LZ��҆�;�1NQF~/�aXfh]�U#��V��9(~����+� �Q{TL�`;�h� ��|c�����C��|���-,�g�W�lת�ND	� vR��%� #�$�O����HL�;`�S�������(�Od��n�2:�"QGލL5��R.!\�o��I����yD�QP1�0x
/y5l����f!6�DH�d֜�/qVm�Ot��~�Oa�{c���MO-9������|���ъ��{r�ݡ�Q\,1��;ZMِ1��'�m�/-Vu=(k�"K��ho��֘A�r`GrD��X��W��#JO��Q\��ꨖ�.p� '����4����DH�����e^ee�D��%:�=��ٿ�}�{��i�'�Y=�~I���H/6�a� ��f���<���<��(����|��z�-C�j�;B3ے�a��w���c�����_������·gQ��8o	�tߌĈ�d	�����q��3a�2�Vt���fM��Ow�!��_J���i4+���S9�.��~��x/x2`�P�j�֝�:A����G���H�We<���a�"l��5�-��\#4��l^Ԫm2B�/�u�ޅ'%��۪�k���r��w�S����қ��c0�]���$�KC�/T?�s��	�J����_�CC�尺�7Z���9�Z�S#$[���xb8�<ź+u���|��.��O��4��ߤT��L�I�0�匷�gJUC��#.|�GNE�a��QW9���(=g_��M����k�Y� N�Jó���Kn�S :A��%�"#9B 
��@�=���Z ��GL�6҉�u�����r!�M��" L({�@�)�hAz�w�$ \�N���l?˽��?O~���4����Z�s�׀�eӶEҸ�SY�>��"gG�۷r�$�����SG�};e%���n����ǂC|VB\2r*���˵�#,HknP��@�Rl�#�#����䧶gXv'��1���hH��,a g�CT������|,ò�P!�xC2"/.�G"�ܿZ��q _��i�����'���8bsr{�"Zv4��Cz��Q;���"1�=����,�]O\?�u$�aL��8�� ><3@�<9�b?�z��ъ����2#��r��}|,+���}$+��ǦZg���0��������`���h�ql�S"#����EWt@�����\��.X������j$-��\�d_���Z��ch
��9�#I$�PJ躨���}�@�*��ϗ����zL�P}:7�>tvC��Ur09�eg_3Q1� uw_�f?;�jT�� ��dP� ����n�Ϸ>(6n#+��Lx�Aۨ-OBl��$8����c;.pt��d�#K��wB�OM�%u�y���)��^;�u@�^%z�`k�I�xJ�Icϗ)���v?���R�k���� 5��C���Q�dP�p�!�V�F�֗^�mN� F� �C�ȣ�di��ҳE�:s��Σ�!���Y`W}��[DCԊ��X��Y��[���ׯdfJ���7���]��W��H�����4�N�����D���뵺ld�Wڡܒ>g�ŇL�U�(?`G�C������:g�{D�N���g�^�^��)f(�lCh���&��'�1��yZ��N9(UPu6#�sx�yd�:����~E��!��F��������#��J��]�;V^R�;(vY�FI~D�VdY�<����mχ�9e+�T�C`K7�O��0B��	v.OŒ2�!���Ϣ9�TP�**L �}ؒ�𺲞N��1�'-ٴL�S��n]��7�:��� g'_����H;+��9GK���b�\��V?6�"���nBzd��a��`�����2���U�6���?/eS`\HU�*�9��"!�����Z�>U2�c�0�^���8�`�RI�#�8s����7"�S1���G��֔�g/fBV�ٜ�Ɋ��'��ҳ�Y��!I?`J5(�/�5����f���0~ELC�ZW���[
-���
�fP4K�[%$���8��)�K(������dޏީ*�ԃ�myC��A@��:cn�}�@�)ev%G�h�Se,��(�пʋhL� ��N_J��P<�7F��Z	\qΞ�848PK��uM�MΦ
:@�~ۍxC�4�����p܉�\Zۙt%���xL���	I)�Qq��,��,Pz��(��5+ؼR�9}��fz����-X�7w'�g!������ �# 9�#����07��N�,�3��[
�lVQ\r��Kݕ��vML9��O{�]E=yyD�G�`�n9�A�/��Wv�2"&(�w�� ��tJ�81���|��H��O�I��<�6�[݇f3t���_Y������dKH/���
2!Q-Y��_���I~7�1�ǒ7)"?��=�2����	�E�W���� ["gc.ޫg����&��BĠ>:mhVKvO4�ݰgN��&�;�l�yAk=�Jn���I�
�ӯ�W�xSM�#�X�l<���
T e���װ�Ae���w�����"x_Ƕ��)�0��3�͍ab@�V�Ŭx�F.��:Ģz�%�/�<�Q�3]�q�:�~7p����2��� �kŠE����U}�?ٷq��RN�F�ڱyN�9�pn4�����Ԉ_&LN)��a=�<65&�*j����Ͽ/)&��&�CA��X�#����YGh�8:j4kD��L�X�x�`<Β�*8
�}ud�5�pD��JrH�B�4K����11�>�,��Qɶ�ԇ�"��/��R5$��)pJ)� J�W���~G'; ��g��Н4���̌�*�� �Z)�1���r)�XݫZH��?>�����\۽�q9f����Q}@��tCu�j$G
X����ac{���!df�$����؇~V���%%�\��Nvs'"���~�
��ֶ�*�/=7)�ڷT��!ѷٳʫ��\��4�O�gI�`��D�P�M��Bt�vlms5�L֚Ʉɸ�ѓ{�_PV����K7�c�pGR袑T f���.����;�Ab��ƭ���iT���%�e�xQB�%�1��v}��R��?k�K��<�K,��"Q��j�	x���0�D��U��|7P���0l���_E&�c����j�5�.�H�a����eW~:�F]����и*ĕ:Z���u�7��˴��	�����,��U���H��`�W'�K#�K�r��-H��j'a$�0�%&p杖a��->�����,�p����4vܵ'G)�����c����kY���T�=�LW��.�}٘�m������g��/r�-eN5k�j͋��R�>w˞3���2��	x({�վd�^�Ud�z��E��4�Sb�R8��Ͷǔq�%��#WX8c6�(�m�8`ɲQ$�W���z�U�w}�����[�� 6pH/Q��KY2w��V���&g;������W
<$gV���\>w|1�H%�[pn���-QJ�=u��J&��:D�5���cw�C���xOb�&;�i�w3��,0��y�c�æ5�oI������8AI����?��r�y�	��uAju#��4���32�X����]Cǃ�.�)Ƃz@�nÊ����������=t{���G�Ѭ5�dBz>[@���<��Yj͍�����t�s}�s��n�8 �D�B��^kr����!��٢e���:l}���_��q�=�Wb���M^�+Zw:�<)K��b���{Z9n޳�J,D�5Ud�*<hE�A*�E(n~^�A�%�<Ό�+�EK��� +���m��6˞ܻ�l�����g�-������p�-�?%G96M�,��M����B����/�GD����_�2n�G��Z�@3����l e�����p���;����/��0�7���e���TE�M|q�WQL;�!�lk�����2̣����BF=>�Y�<?q����r��Rjy���e��0�C�}ȢN<���;.ݍxn�[ɣ:�9l5e�6����]T�2��7��r�ɔ?�p�|� ���qMoQ����@��,8�.k�NieP�&�f����
�Ur�����ML�	�@�
�Ty�
eד݁�|`�9c^]ڂ�H1=F�H��坤��b:p[��oZ��_x�s�yv"2Λ��1maC_�oҍ��isT�@�6f�H��7�v�>B��n�A��[ғ��fݥ�s�P��u#�m��z���*�����SE��j>�X��oY��Eg��K���.K�G�/o��B/X��X��+]���@�����EZu�]����ܱ�%U�h�B�}���.սD.'���k'��z�k#���{!���~;��N��~��'iںf�ӆ���i������Ѿ6�N��q�571�NR�k�J�ݞ�`<޴������|o��=�zFh�����">��"8�A���ы����q�
���r���*��l|�k!�Xkzn�4�0*���=��h	As>���/#������`�v2��n~�2���[�q����`��E�{f��&���#f��u8_XQ��v�'�p����ieu��g>�
0����+CS�; ����L�>��r�=FīB����LB��>[�^,T�Ѝ	�����r��.�h%ٛKl$�1�ƀ�U����j�M �Tfǉ�o������ooc3k�"�q����v��M�n�wC�I�Br ��#OFP��N;�1�����y笵��έ-aI2U���+���D��ۓ�Z�X�����F�S�:!
�eM'�cj��dD��Q�30x�̃+���!zf4 �H���*�*����4�ʗ����4�A'd������
�T���c絝,�j,b����d���|��N��8�DY�=d����L���!�٥A��t�@a��W�sm�{��+y��֚~��`�B�K��n�-�Q(�0	_MG����Z@��~�B?=�t��b���ܙS�
UI�il?bº����GZ�n�W8����"T^Ԩ 2���(R,� bj|L���)Dվ{yj�Re�w�@2=�3p��h�Əii0نA�W�V��	z����.CAȸ�y,���B�1G[��&���N tl���qh/����;I�sOp,�zJB�Xt^�ND���i�� ����^�P�>�F��(�$[qًc��B���h�p�89.؉��{�����o�ݦ�#����t�)^!}����M�Yff{YMe���'I��w`��ïh���H}����M��	��������'-U���6�-�^NsEK�>����]��%�� c����&�'ݰ�.T�C�l���n���`:������>C�v�P������#�&�<�1ފ�R��Ɖ"�AD5ܡ=��m�J�E���_�z�pN�}�G"��P�쳹������H�����xx�x�MJnc-���c�NK)�M(j����;�|�#�Eչ�,�c�ZS�����8K���(>I���H9�nv��e�P�x��k*M�cvʐ2��դ�dJ[��U
���5	�a}�~�C�#,sd����]�/b_k���8���� Ah�
])�v�8#"N�e��2��m��x�1t�<	v4��$d���R^Jy ��X3���|Yr�/L�\UA�faG�$�����fe��°?[sz�I�G&���rU������A⫤��F�=V�R�q���<ń�q�	q�#邗�o_��B�.f_�c�
F���Fή����nIAЅ��M_��G���A���@\m����64��Q��i�k�{��1�T���Z(��q�Z�4�FL�ʙwÉ۟	ެ#e�"f�g�\ހ�z�{H3Xu�w�꾿�R=b�#����� S�1Q
VH)'�h��ԩ�.|�J_����щ�N��ü�;��X��B�����S�˝��m��$j/�-"a�B��r���׾Z;خE�XҀ�9tp�O
̡�7��m�x���,�p�r���.�7���p�����&�C���1@�YoV�~"lz.�)�{�#�^�K�.��"��x���`�O���'3�.ݗ �/\���~%1lm2�QZ�j�Q�2�}�ߘ�4���� Z��I�My��
�h�=֯�c���#&��ړ��0����;*�ΰ��������h��(K�l��Z�xۃ�w�A��O����\PI�EM�r']\^	#)����݇Z ܊M>AR�*����+��x��P[*�]������Vu<�tc������¢Ϧ�|/`�R.吿�"����'�{vy�k�B(���3?�n#:~7�q_�͐�8L���E+������� �	<�^�p�'��eɦf�6�ˤ����|]�����u:i��8��G��t�^��-��m�U�������G�F�:��M�������
��{JzUXZ��ba��6�$B�`�+=M��}�g��- h�k8�x}�4��]Tg���C�H�49I��>�ԧ ����5���(t������꽇I>vbz�n��Q�2��+r%���me�;���Z�<	�ר�㮋��泽���؟-�'k��z'xp�)ޓg������^ʊl�t��(�w�/A���u�\;�r��\��)����Z�~�X��xi�p-��S���)~Q0��b� �zl���[�wGB���c�����#��H?��k|�޺�!1�x��@/�&�����7�mwUi�ƠY:#ۦZ�#������Q cȪMxǚl|2f����˩Q}���@rx_ߨ����x9J�r���)���L��u]Y�L�S֌���f�L���.��v���v�J��ٓ]��J�j�.t���T@	��'��
��$o�=�R� 5ո��y��7�oݳ�jjy�s78���W�Ʌ�!�0a��r��C��F���@V�OmkHr�ub�%��+�5�@�gve������&�2�~���u4�`0�˳*��3�a�R�kd��4�P�(�P���[��\X�!�� �� E��E��;�d[�Sl�|��=�_�	q����~�<8	��s7t��v)��#�L�����%���1}5�"L)�Ƶ8_vsaۀ�F;�>�� =W�э�޴�ʋ.����p�I����gKb	��z\tY�j�;���H��5Jw(M�Yy���&���lA�N��5���YZ�ǡ�$�Y��	-x<��®�PQ����NSo���Eһu��+�0?�i��P�^���HKU���pD�ar昜�os)�Õ��i��U����O���A�H!�K4j�35�*�w����xҠ73)^B�zn=�G��������>T���K0=�&���$qh�5e���̽h�-՛�?�pk|ߨ�8���,�s�*Uh�'���_��g��ٓ�1��>3�^�D��"a���Ǝ����H�9X4���.CFj�#.*�R[d�q���S���kx����������J�T�b��<��fY1���!��Ƒ�q��n2�o�=`K��>���'���?٘0����_�8�>��0��	�7�y'x��$�c���[�ڰ"R:{x_X��V%L`��_#�t�1ќb�q���FТ�gL!��)��P!P:������<}g����_��a�ֆ8m.n��[!�1$b��c\��jg��~���Dk��/��g�%�L���3��-\�TI3~�����<!�Y6�|�J|���QϬl)�l|ۈ-�A`!�ql��%!8j?��̈�@�a�	"6����e�{l��۷M���).��y�qv�{�8�(�b �&a�����������|v*�z�D�=cY�"�����T��U�!C�	h4��4>�ܓ�9$��Oju���3��~�D��؃�Bw��$Y�ݵJ�Q�b-ߊ[�}�`wl�%j��BE%�]�:����=,�s�ϭA7�]�8fό�aJ�	��֙�c�mt��vՅg���>Y��k�}�vP{�5V��;���1������x�d�t.�-���6�Z�\�A�׬�
)'�7Y�̖�O��������^�Ys���-̲���ǡ�H]���/XO�*E���l�.(*�};�3�9Z?�!���L�D1�phv�m�4n�Q�yl�k%!��{�'8�5��Z��5g�����^:�{up�w��n>p$8 
i/?���~X��U��b�M��>��#����>ġ�H���Th�Wq�����w:��\h�ڄp�Za�o��������]�	8shJ�T֥��@�:��Q}f����v�U[[�Ԡ�������/���u3�I}v��Iw�y����-� �'ͼ+2��ؽ�ה	��l���]:</��}�n���/�|�4�I�b�g��яߙq@=��˯x6�����]���\V�}o�"��ӥ�	W��ӯo4F�>h�s��r"=�8_O%MbE�h�^E��4l��Ev$|���>�>��ֳ�q�2�����rG]-Q�&��Xޡk�G�6�4S:��[V�L�K�����Z{�y��-W�8����$�yp�vˆ_;nٿ*���Z�=2���K�N���X-��>����k6�/U��{t�= ##Ȫ��Tn��u��NP�}
G/%j{��Fx����ǉ{��e��.��q)��"�@B����R(����=���F�K�r���A�ɜV��I=�W�υ��奛�AA�͑a|�p���I;�]Z+h}�c3*|�E V��3G3�R?��#�#W'*�)Od�<'��UI���*?�:$�c��Xt��c���>�@fJ6�|��9����)����Q�x��ua[�� �:{ms�μR��z��y�&��Zp��Ǝ����B�9
����n��Ϛ��{�Ҭ��Q��C_�m�?<b�^`����Č�}?��)�}��f$%`H�cw�\��1M�%e-��}m�2��c|�ׁa��̉���I^���v���s�H���@�Z���\#�«c��XF}�i�Q��Y�`sl[u�� H'B^�-�f�@�R�WU����( @s���)NSϲ��s��2��=��Ȏ��6�n�[�_s6/���2C໿����>�:W���C�w��#������,,�ϴN�� ⑌�-E�Z-��Ŵ�����;��5�:�ԑC�*�f�F��)���@�Q���mn��&��Q�:A.�
�j9o(��Rc[��;ә$ϧ%T�� ��l�F�>K��0.6yX�ϕp}�	�Ut�"�(b��[�#V3* ��e�R��V(�&���.�"�=�.3
�j(�L��Um�c..-M��>Ew�?	��3d��x=~pP%�Rp���cܵʄ]&/D	.��e?Ny�U�V�y6Y��ʡv��/iZ�	�#G)Ȭ��@�M����CQ��d�_�\�EU���1�� ��X,M�X�%tF
5S��U��+�E��Xq�-��]��_�%��*.
�(
�<�T�`裮E)`���v��(�g���0=-�p�6Qw�MJ�/GE3 j#v�Ӟ�[<�^�>(D�*��!6�.F�$L |ç�6qɋG��5N$lH�V+yZ�53!P	o�,;4&�,��^.�����.��\nD�:�d��H���6�?1�ű��m~AO0�6iT�@!2˅��hz�aO�²*�1��Obœx+��ְ��>�|�̠��`��>ނ5����^�2�,����?�r���4�w.�
 ��`�lb���`��A�m8�:>5 �I�RV�({��upħ	�%s&��_���P��X�>�i-�
��Z*(?�eVo��\U����o跚ܳA��L�N}��'7�e�j�9��'���oWxn���e�P����)���Z�ǁ�;{%-(���A]��k���%�"��n׹�����i��·9����*��b+�Jr��L�%��T��k!��9g"B�ުJ�e���m7�s>��IC��C��݉��o8�w�²A,�ȜU[\��|;���^��X��79PFDaѝ���o�Z|�Y�e4����R�Qp����H�S�j%����,�i�0��k9D�r�F���u�����U�M+������G�� !��k_� ��H�K5)�FPz	W��o�ّo��d�����Q���q@6?W�<��'��[(���h��}�/Y�{"͚�q�WF.�$���b���X��k}��Ze�:�%d�z�d�`�X��o�����UɻZ�k�c��3/��o?�
ņ	���Z
��کMz�I$��/Jk��h�#�j��z)x�?h���D(X\���U��Rab�f8u<�o���-=�Z"��@sW-����Z���.��j�����|�/G����F��
��V|R�&0����o��>X��wugSV�rS:�sU-�ź�`��2�.��cx#�҈~>�;������CumM��p�J_�ܕN�;J ��}W��(2����ۡ��NV��P)2@5���E��ľ�ɰ_#β"_t��h[f�[u�O�a^7��@4�L�Iwl{����BRDW���G��q-U�5j{c���6����\&@�&մ�5��ʹa��{z��!��sM]L�-��Ҟ/C'������,W��=�|�ʔ���]��\�F{QL�u��D��!e��W,��=�r��b���*��<�{���?�
��ͷG����s��)��%��:���Z�}�6��N?>�1��R��PU}f5�]�Z��o+�� ����=奷�.ݩ�%��`���]��l� �똘�����/^(����v���%�ȕ8�/ϝEu&C��o/w��5V�!��!{������!��O��e.�qZ���R���/��`���b��� l4�2cH�usif ad���s�>�v?�nG`)̝���a�w��?���C�ۻTk"�,��=+l��R
��+ΒQ�����q)&�q�x6lf��{�BK����!HWW�|�1 �,�����' +�;�j�S�eǝ�]����NݑI�#o&J��ٻ�B\����"#�8��:��&��r����-ū�y}��⦻�`��q��4�`6�f�O������U��˃7E�`�΃��2[A��Q+�(�t�T�LC(���l�Z�+K��&��4E�t�-��e�9��T9�6����r0b�˰�s��3ǈ���Ɵ��������S�8>�>q�z���w����2A
vȳ4�fqd�RF�%��x��T{'dЅ�kg�*;��oz�=֐���~�)�:��K����i��FwWd~�O��A�a	u�u�N��ҳ�"ɥ�y�4�R�A�PY�P{:��˚ٜM�چ��9��~xM���bAig6���h��<z|kw�Ņ��a���(�|��wn���˨"��/5$Kn�*|:���f��	�'�ȧ��P:��!�@
���0�Ann'��8ByI�w=.�f4l�V�8���G��x7s�qoe�@6�dpò`��-r�����(xQ�Ai`���i�{yFI�hl����\f��c��ŋ�V�����@I½C�χa8�R�� �_BI�ݰ�y)�D��+�r3�	6�
���^���#���w/*���-�����Gwc�YJ�3{���1��!6?KO!ɗ�o����@�?��[K5/��i����|���^��Ժ�]�/ai���n�����*�t���J#�S1�y&=JT��w�wӉ�J�AO���%�����ypq��c��O��v�s<�),��\X4Z8��k֧��]O!W1t��04�f�P�r;q�������V"Oy�^M����sw����ڭ�$����Z���	�+�h�pߥ���[�I�9�����3�_Çi����h�sͺF�'��E��W���9=IeB�����c�nv�e�&�ʐ�z�i���o˗�	?sR�ŏPɞ�q�;y�\�E���mM��H�r��z�6���2�!d�T͟pౢ{�;W�{�+	]%ˁ�8��{Q�0[r�<�����!��{�����3�������U��\QA�B:�a/�J�7�����G����V$x�Q��O�}0�,����ZG��xW�G��`.�{�g��=�	�A��vJ'�J����k�)~vz u|Z��}�1��WN��F�SJ�	#Apeȴ�:x�'|e��Qߒ�u,Y��Tn}G�4�>Ł.u�88vJ�Y�v���,�n������%[��,�S����A�%G����5U�0���K���_�(��ɭh�۩y;mɤ�
�I@ -�{l�]��Ά]��JxH=d�&�牃q}�윕����� f�R7���4�_�.�n��|�-|�d���O�O,1�.4J�!�Fƥ��-��NX=�ͷ؜�eL��W���f?��Ŕ1�n�̦��=:2V�����7[��l�ʁ�8#R�w�Hm
fT�������,]�Q(��c?���u������R�~��#|�l$��L���}6����C��]g��7�Q) �{Hrs��������È�" R��Sk_1�BU�1H ��=��`�zB�����frю#�Tz������	Q�q��%�s�cO�R<�G�ô.s-��v?d���������_��_Hx���.��f�\�<�čJ�2D����>X�$�9�X^�	�]`B><�H(����~i%uM����J���'��˾WRSGP�~hS�-ID=T�7�9ܗ��H��WA�}YHZF��/9��L>�m1�Y1���;1���4H9�a��v���*:��B=E��0B�#w�Rj�k|�,CQ�1���K��Ql�)��ށ��	l�:�׀
9�"F��������q0g]b��g�������}�H�����݂/gDy_�i?��׏S�~�(���������\0������r�\�������bl C��4B�����5�"2�;�S��UCU~�̚E��Q���^��<�(y��hg��{fqL���f�7b�B�t�t��2��)�ZB����֙4;߶C��E+�=8����c�o�ы�\7�����lv��w�%?��Ɲ񤑸V�+`�	���	K4ŻF����6� E��u���W�D:z��V���4ܩ.,�3��9��O�a��!k���jR�|Ϊ6"Eű�4R;ai�%��Ư�h����=C��7q�����%�h���J%���U����b+ �2�K�75Kn�"��Y?�Y�L%Hn��T�B�vn�2�f
FC��H�DZ_��j�����e�3	��~�S�h,PȎ����q[pb��M�dN�G#�5��hw B��4H.]��D;i<�����2����;����wj��_�a�\�7&%���N��B�ʢ��~�c�K��൳R��U��,e����h����p3;����m|������Q�CkO�JY���n�^�����NH�~���4S&ԯbn����)֦\�-'��*L��i�m@����T⍓y� �P¸&9T�n[�D'���bkq��z��ʿ���l,X���
|@s����!mߪ*M��CY���ؐ���� �]2�*�ξ�e��ίL�Pmf�!H��f=�E��u���4�뽄�>�1�o��c1���Y.zq�R܉k�50cGU��[�ʈ���$�yC��E�y_��ď�#,��\"�Y#� {V��m�{����dW 1���*<��؀x��Ζ.j����f�A;FF/rii��?+�QrV�5>x�#17s��6���lZ�ȥ7ݷk]d���Tr��?�⒭���A��������2�2��8�\F��RaQ"��qR����;/ݙ�^ؕ[峐lX����Pc�ԭʦQ=6M$��E>�t�yr�sBC�i(a�z���_>/p�'�s�N��@��\�2Y�2�ݱM��Zx	���*6��{�@�~V�8���J~lv��Equs�#��Qh��c�J�)���@�<u'�#��<��'���7H���s��zK���a��<Ű�h�v5��s�W��������5�u��1?������&�J����|,�K4p�Hr�bTS.Փ������ ~����b�����/��o�z]M�_k�U+~�=$�&��@���6��?�5A`���+��*)%�p�g�[�kv�vS���l�SJ��&�YL�8�1C	�o�cd��vyP�Q���}�ũ�[���<=t�D��g@��� M�o$�aB�*���ۚ���S9�~�����p�G�M�`A4�-
ޫ���f��pQ������>=SQ��)�K�P�+��#�M�na6I���אd�h	��Z�c�@�)�OE����O ��N�s�i�4H��#X-�(K���k&gsh��j��������1��\�`��a���f��l��c�?޽B���Z���R���3&S������f��ژ����`YDOol���2��9QT�pi	߈D�i$�T�/i	I۟}�@"����.��sV�-t��F%,��ۆxr�� ;�ŝ���\�&!^w�Z��&u����D��>��:~��'.��L�9�Bd�W�,�[ˬ,�닠̘r���U������#���C!1�ds��g@�n��:i�-�p4nBVXd�P�nB�������v]��%e�s���S�m��~CAg�N��r�`t(f��ÝQ  7/��YK^��7SbaO��r��[(&��5t[�����!���R$�ȳ7���=ԼrQ?bFkGC�N�����7��=��I���H�U/L?����gN���~��B�� ����v���?6�$l�5�9UV���K���!yb|k��!N^&���o7�B�Vȍ��	�\gG� 	: �D;��]囶
!
��y�5_9Kkh@1,���z��!�uM3K�G���A���3_HOD�P�%�g����1�c��a�����T�n�v��V�%��YSd5x��ො�{�<�Zj�Yx$6)�*%����yN1(/a��B 8�3(y]x��_ 0?�-H��U9|�xg!L���d���uk����L�{�?͐�*�K�h*W��������}�����r�E_��RF��ot���D{�-�1<[4O�1��/���#��y﹕���	eD��/����t*V!tK�=b�YP�$YRx���+]^���wrDU��J�a��b��]����!�܃3���&��tV�O�ݯ�P����i~��t�:l#pm *�AJ� �w#��u 7� y\������E��ƌQ	�D�8ޏ��.���)���υ3�[�j��u;�X ('����R��P�}�p��)���.�;9�WH>fERJ�(l�j԰aѧ��8L�mN���xE��IP�d"=��2k �5�p5$ߢ���)u+�­�`�/<	��~i���B�vl�T�W��֥{�;�
z��9T���J� W_�$k.ݝ~���!�v
��p��@�KH�U�/��	�Ȫ��Z��=[����#z�"?o���s�𿤜,��$����Vj�����"=�;��֜��g\�Y����/r�X�B��yC���ʡ�K���:�/!'�&ہ`��s6��O�P�L�day%r�AM�~�w�����B�3��i�V�蕵��Sն�д�tnT1.!��i=����lM����4���Qh��[P�+#�M/8�m�����#G$�X�1U�W��b�3z*�ʔ0�6��m��շX��~��g�W�xaVB��L.�Ⱦ�#�#��n��G�$UK\x�1Ԅ���Т���H�/Y��/��j�\ �D��:ꩾ?n޿��Q3���;�-��I
�*��\��w�᲏��c��ѓq��"���L�"v���uqw!�	�!h�H�u��ȉ޷'<m*����r��QH|m�<N$��8n��ƣ���A�l@p��.�ܼGhH���6Dǟ�j��f�q��ż|��h�Z��d,���<w�٩�'�#N?��Y���d3i�h���!4K����205���vD�p�ٗ�Qi
-hŊ$��ymN�3�Ъ�ad�ts-�!�-0yX���9�-a'q�p����5����y�2�W��P�7�&�$�Zh����,�df_��Fq�A�&�����^���v~�z뀆��$΂n0�0�|�.|����	z{�(�7kP`c2�Z�Feًi�u7긴8�=Μ0�^f�>��t��놄��Q0���ĭ�P��}+M؅I�\-W�P
T�]��a���.��h��??�+U8���#��jK����i��k:��a��Z��e�ɀCLT���U(��`8�Ë�?`���B�I�\|s|�)ϥ^]�m�4M����{C���>w�'2{��o�U���`�f>J����������d�9� �G�Sa�ڳ��tDYv�!+��2n��By���=؝�C��+>�;#�s�v�B�
t̀���{1��'g�t�j̝�*�b�$��դ�_���T�k���衜G��E�H+MUa�a
���>4p�WU2���<
�{$��'�':6/�5�Ds�c������_
�͗IP�<若Y�B8�L�oz���%M��1s"��0BGנPP�۶�n�s�'��X��b�����e��qi��"��E7-4mnE ��s�_��0��v%F��M.-K^
�Z����ØM`e�Z�ȩ�_Ѣ��:m'�vD�]֣eƛ�W�#B��N4�R�{څ�Js�k��ډ�>đ�a�S�m;q
�1�R/�(�o!Z#�,.�N2�hw�wy�)V�gYN(g�����޲f�i	+�(��a�S����3����_�q�+7s�+�o��"�:��bG�yR��N��x<C	k����JURE-iUM�Is��ʁ��"4�H?��ʴ���k�d8�ov��J��l�%�h�9��ޕ}un�4���=����2n�\y�O���\p5��]����+םeIsX��7�0���'���X�kr�f�'jNٗ�q�9+����zÕ���ChFt����}�s��������TQa�P�p>\h����F�y����CT8&0�:F\Ӌ��<
�W�ya<�����H�gF.x�f
y�;�uc�����B����^��L�����Oc9K~9zb��N��5�|�ն��M��u,||f\�yH/���b���]C�����p��E;3a��
����+Bc�*-�j�����bݬ���c4�03�����wK��Tj��@l9&��'uv�kfM3���zs���K�FVB���0����anK�0B��K�\��+�/�����Jt�k�	k<��q=>Y���F�u���G�)[*F��[���E�0�-d���(�fJU�%l�<C�["�ҡ���\͸��9ޓk�tή��clŬ�Vd�ԮΫ�8����n�o#��5���D����{	�P��m(	�����(5eb����M����ͼ�������@&�7�(EnWR������/�j~9 ��ew�B�|)$���!��H̳c�e�G�� �������
&�U�0���*�$ǚ��������L��0�ќ8��_�RO��;|8�/���N�7��%�&hƳ����&�Hn��l�<�Ȅ�p���2��L�}�_ecs�P�Hu�*�,�R]����DA ���3&��R��s1D����xx��hp��OS�3�4���}jA*4^��`��K���ۏF������K��h�o*L':,���x���$�4s�?���4�tUD�H&�8H�_�Z�X�na$����WI�#��a��{�U�zy�d@�N2֏�"�X}���z-K}����L��HR����C�]��Ԡ��c�lEs%0�q�n�K������.�1g���}��=����
����s8(�F�w������})\�'��B��KN��8"��v �o����m�y��"�U�.%T�5`��h7�_�[�i�i�fv��Y��k4G ���$8>�* �����v6��L�+O�>TM��{��@ ���P� ��E�*S������1���@��?��֟�@Hy0C��{�&ꔽȁm*����%�?C��e�D���U4d&�|��+}��8���'&�����-vZ5��s}�=�i^}mR!�
��Q�-��{ˬ\�ޔx��[ž��<4�<�b�\�t�{��$�Q�^%Qǧ����I_��
|x��4u�P*��9D�)s5��D����k�+i�ud,\�1S�^����6�#��1�9ؒ�*�W:
�0Er��!�wS�K���S�&#`Ԯ]����P]{����c����F�|2���\�.M�F\��V�f�$c�2����v���(M�
SA,�;�"��I��D��,��\j�B������ݧ�?����C���f�@�Ἂ4�6�9�B��K��S`!�S-�e��Hc��Q��4ϫ$6�y�E�)�������&2��<�ͯY��m��P4u#H	2E�G�}����OTC.d׎�v��9��B�F�h�I�3$�W	(hD�2�Jg	il[�����&��������ӂ�~>���܋�r�Cca���R�X������B�'�:����:j}dWB �;j��Q�f|:���@M�2�T�n��8[�|�~�p��*�]�S�>pP�\1�K�5;̱�怺����hv���_4���k����|`�,žw�b�\�K/j��;���ַ��ַdZY4CkZ�Iw*�������:p���_�R'�	O�y��<�|��$���b9J�f�Zk� �#r�~�t��< ����	Ώ����EE���w�{��[��>7�d:j���g�����=[�!d��Q�YB�.��:��/,&!���^���S�Z��=�xޏ
�DR���7���Ib������Xb�X�����D�y�'
"Y��b4�&v�y���'o��T�ĵ���h/![�
�εeݒ-`6��n��T��8e��� m���-�`��W�j>����AU�S_���.��9) �sN��ZS��Q����w�����tR��Z�:�\�xĝX���6}t!�i2)�J�ʵ���gE�����	���KK�s�1 _���'Wɹ�}A�Hc�1Py�ֽ꣰=�Bު'�����o���d��̾���3ж��$0����kc�wuS�DY���S�/�h�C|p.6ɓl��1?�vN�[S���>ce��w��\��?g��/�EM�5�=���`p�M���
�D&�s��͋�����IVS���[�II��D�wR�cf�
�#��u�$9��z��MHgZ�	�R�M�s86��FF�1��m���&k�n����˗k���(q���I���a�\���G�cB�����<�j���L�P�V���ŏ���^~��u
��W)�;NSt���RUW��d �5��-%!��eH�9w�q�iS.K���N��P�0����!�Y����?T0P �D�},����%&��}�B s�y]tK5��/���zZ��2�q��ς���(�7��
;�b��raS��O�3X+�l>��u�zn��9ʏr�������t�-� ҏ���k��6_W�2 ��@�Ђ�{����N;���"��0R��*h�o`�a��	��u���1�a*;Т���ᔪ�Ƭ�4[m*��R��
^�3� �脘���|<�O���Q@�o�(M�5���H��3���6�������,>��+t+�H���iG+6lvT���ޢ�zEI]��?��֙Q�H�U�nf�冏�!�=�E�{,`��P�"�B�FP�;}�O����o��=MpC̝vh� >Ix��Q��Y+e��ǴL~|`��g�|(��[��A�����5k��7�`,��[�Z�����Tҫ�H\�}���}u 9@g(��؈�x��j� ��b�(��.���V�Z��&ܜۀ��o�����W�۽��C;�l����6SOQl�`Sm�ck�֜����h�c�t���Fq@�W���N�$k��-�H������ђ�&��?��$�8J}����`,�`��T���#�Q,6�l�u1���f0�~�	�X��뀿6YE�=%���ת��mtc�zPf ��d�5$��\]4�H+��>Y>x�/�_L�'�,�R$p���N�h�	����g@Z��̂,VۚQ
�.iK�������$�C������aY��%*q�^�}��d���B�w�:�NgV��ED��9�1����,Hx��n��ե�p"�^B0lcPm�z��ɷCH�)�Ϩ访J���#L�d����R��?�ys�*|��^.�/Ƣ���9_������H�ޚ��q�pN;�+��o���]v�N�Z��tmN���R������*����֘�C%��̳Vq�T�.�ܬ�[[i	��h,�&Yh|�6��{M�����g�SBuՑ�����7�vtm+[�~&���~�
N�(��l�a��fA��8fb�2�Q��_-K�+�Z	�l���<ȷ��cIw����7@g�,�K�'���Y]�I�"3��d���.p�w��s��8PT�r"7o��`^
�r��J%��BA��/�/�	�7S3��'��Y���a�=zj�]�w1#E�W�Qý/ܮ	�8$�i�
�9$CzC�r� >�TR�&=�]4^�E_�>����jټ�?S��L|�*!�9�\GS��E"N(4��x�A���� ���b\,k!��M��;N�3z����uT��G��:?&����3Nҡ������o�T]��Q�]�xa�Ȗ�cԟ>�����`.҆	jޕCF���3A�U瀯sؓ�Bs)Dg�r/�MB! N5��>}��~��Zn�&|S��/?4�3�xLa}[�<i�S�=V�Vv(���A^]�1v}�h.��'�nL�ѶJ���(��:�_@��m�L�?YX�ӽ��՛�����>'�N;:UJ*%2sz9"���G���_m�':/�&�����Y�jQfU)���t�)��YS��D�>~
�p�V\��W��A�,��+�W*_n���ð�!�l�z[5a�� ������=��p��Wn���Ύ�p��oMP=�=�r�^���v/�v�8ú�8��l �V�ƾ%@�`��8ky�'vk����>�h�%Z�n��#i #��Q�k��Ui�Y�2�_i�;�A�^[5*�׷�\��^=�n4騢��{�!a3�Ơ5X
�$ULE��(-)E�lEz�ӓQ��C��#�æ��5��٧���Qİ�T/8L�V�y/Qwu�����*��'�~c�	Z�8�� !'C%7��_�鶴�j�rM;	�aX'�z�U��ǌ��X
A��3V%�q��nNx�Ếb��[GC��;��L�r�GT���n�r�8�Ǿ��2��y�4�$W����y�"\�����E\�EF��w�J��CG&����-
�B��P��r�
;LDYA� ����:D@v��p����/��O��ǣD������:��<T���z���x�)!:�ۗ���ŕ��?~��@w7��gʑY��.�]y��gM�u�^gJ:s�[=
����g�Kz�X�p��4���3�<������u/=3��� ������CQ��Ehv�_�:�{�U����Ae>��G�OxT=o��:r﹕�B��ʴ<��*���%��?g�ݳS���	��)� ����&G���r�z�Х���a��j�Aձ��џ��ެMs����Hy�g�ຨ�]���7Oaf]�}YP���x�����	��ڲ'������F��px�t�w4�Nd*��<��M��XUU��߬ DGљ��K���:�#%�k�Md�]
t���.~[��b$�c˛�
�uEL
	@��ݝ� J`�,Q��Q"Y��M_�l�NA���[F})���gA@��/��� ��Qϗ�!	�Z^���Ot���@���鄣q�K��-n^~���Y	�"��91������ӭ�X�;'7S�r�čd��7��ǿ5�ܒt�ہc���j`�c�ng�Z�=�����N�{��� $��%��YU���%��؞�Ӂt���5;[�} �'C�w��ύ�/Oݥ�����}}j2��XYf�*�7ɍ�'Kz���,���lP���:�֚ 5O$�KXF�#��a%�p��*�Yߺ��w0�:���U��#W /�9헥ƺ��������_���u�W^�utZ�"E`�ђ�Ԗ�'m����V���ň���v���<��v�n@&�s4a5�2�3�)������2�O�X���qj�Ji'�AT-?�����j;.���{X����9�n%+���b�1Ʌn����]��[�a|��O�"	0j�z �dj�wR�l@>�<ߎ�����9�c)V@�Ai��p  �_�e���)��t��V�u�F�uє�rWE��M�H>2�F�Te��؉��,����'������I�
�et
W~�����nvR�b�7�?�2��у�g_<�p��A񯦽Ɣ�T�x6�O[vU wo�c�[M�Ph���P[[�A��o�ZǻR>�d= E�7����R�w�<��˒�SIrO�rc��:�G]��� �uB����%��2Bn�l�z�A�a���B�Z��؍�]�(�|�Dr^T5K�ﷶ�� j�*���3���ȳ��ʆe�	�U�[݊�3�֬
�"��L�]XۛܜBe"#�$��|<����YJ��D������u�;6oI�Tv�$k�[����GX�ѲI�ܱh��X�p��S�/~r�ib�]����2jٹ�C�C�"�n���T�M?LB%.��j�%�+�q0����e�����D@��I�V��M�Ui�)n�fvnε�W���%Ԏ�7
2̎%���C�n>9�e!��m�K�k��p8'�d����|p��é�:E�^sh��'@�^�pߖ�ϋ% ¬:�;�>s�W�I�?�*��T��a�4�#��N��V�&�6���2�t �=k��ْ��\`l��o��I�C��%�,Q/
A ]��t�P�Mxl�Y
L��!��)G~�P��	@�RE��O�Rχ��^��+j=�p@��7y�Й?vˇ>E�8��e���,��#i��s��u�!�r��ܘY�����Ԗ���ɹ�mFsL�JkH�gʢf٠����J�X�;��h={u�%0q
?��P0���!Vq���r�^ A���|N_�:Q��P�&��mw#�'XC�Α59�6�3??#�	�ݿ���H�Z�O3ǭ*O�3��N��Z�
:�e�e�e��!�__�-2�6��M)�0mW�pbL��(�����*7f�qE�]P@��I��7k��k�����Q���@0%�N�=\T���Z�͆���~�V�gV�`�
,�c����Oޯ!9��N����l���=�U�mS�ܺ��ǼB))dA���W.�������)o"�)ͦ�#*]I= �0H�{������{*l�0�2�I�[�U�7��*I\��X�5�,��']T�!/�\�C��H�!�~PRs��(����Jr�*�HOՍ�x����h��wC����ՉڱL�GZS�7�X���)��g_!;#��Kn�RB��q��D������Z��\('R��M��5>�Q����E(M��{K(A�lzF�ĩ�t>�u2��}��%y\��\E���5�2}qR[vCS��d9K�+k�����*ܶk|���V��4wS��{�����8%���H5
�R�/}9�-�!���Zw<�[Bp��%؍�fQ��p ����)�9x g�~R�]08B #A���k��-t��#N�Ԫ�[�;͠�SO權���װ�Ќ��.C�:(�+��F�c:1�n1��mip�RP��`=�f�������=��ړ�L+��W���]!��o�3�J�K6B��F��O�e'�X��nS�L@��ýiZ�=�|��iS���YP�v��ۻ��5��CË�~0�n���D��WՉ�F��> �MI��1���AK6#
"���=��T�A���c�/�R�J�j>�=�զq��#J�jz���a9����4,�|ࡘ\i!y��^���h4Af�8��<��n'�����L�{��}�dK7�Z�w6Q������ ���o�;�Z1����"��
���#T^�+1�����XB�&��»&L�I�"��Smb��٨߸V�SpTBA�W2�V=PF��j�o�$�fs�Ԭbh�)��6��ޮ�?/�՟S7�CI�����J�����+�ފ(]�l�4B�7j�����6�>��P�Րr$8���M�t3�T���7zM֌U ��`n������͈�Mä*�ޜ<nEۚ�ZYΔh�Zr =%n�>_��r����	�fO���>[�ENC��|�4�]�ُ� �߼����޳��]�����D��W=+���6��#?����|�[^Ԑ�E�V��n͸t2�`	��,�Du@0���o��0ȋn�8���o�� ʏYJ�k`YQ�&@{���؀T*�_�!������2�ė�f>+d��+�����<N���)�Q��H�~r,q���%��*nd�dͨIO��M����04���=g�d{��N+O���ǡ�R�ߪ 2
���p*h��75�w*���s��S��TGxe��Y�	{�]���Z��^'	�e�����y��$:ל���uj{�8c+�����%�6`m�~@��Q�Iqs�7?}��j�[��_$�n��0�W�JUyn�w�p�џ��ɕt^z*D�ߌ�k�N�b��/�U���h�)A�E��7(�N�Kڌc|��6�/�L��YvŢ|�B4Ϟ4{A�Z���S��\��L�����x�k
������9#.H;`��IN&H���F����R�b}^�ya_M|��E[�~�{D�~�yAN��7������-#ȿoې�t�~��l�.jm�p�6���zRDh����"a�n(X˧`�S�]bQLj����`�fIC��T�C� �T-n�m���$�����SӬ��$#w��$U���ތ�G�]K��N������:H���H���	�z6O6�PoS[gFs��9R_��1\]a1ig.���N��!��S�~�<�+9���)�z�+ �*�t�nS��i�|�<���-ٴ�\=�$���Q�T�}�3��i��g�!��D����<[dL��O��e�1]��9]����(iψtq�����Xz�$�Kٌ�z�ң�oØ8�����g� ;vٛ �q
(��Oow�rsJ��+܋����C�Q��@�/�Y ����<t�$՘�]2dW�ުf��}h)�S_�OQh�z�V�^1�w���ϳW'����1�6�xS��=�$.��oQI��TC/�ݻ��N�c���i�~���&t���ڴ5�[�]��%a�^�`vw}��Hإt�a�Lx�`~���I���/��fp�'Q��:���M>�kMYbi�WJ��a�K����"�;��$s��2�l����睌T�f�	����$A9O�'�z.ڀ	��<6�ٓvL�^��K��u8Hw�76��6�yE�F)��A�ZAO� �Y�s�H`�)������<#D��LW��|d�ђ�t����X��ԇ7�Ϭ}(�2����Wz��[ vv����������������V�x���Q|"� ��,��6���	 �`eN;x�3��% ���˙��dU�:��Uc~��ϤL�C�7Ž�f�(e%�#�R�h�eAa��	޶��t%\�t�-���j�C�"���q���$�v�_٠h��M�%b,2(��	�8"sp�W��2JT+e�]�⼾�:����
����	&Ey���ҿ����㪪G�g"�2���C��v��4L��ǚLY��W�YjɄ��H�,��
�#1�X:G��K2M��&Z�!��1���V��j*e=��x��5y��n�0�ڣ�}�2�+gh�bV+�$dG�a�I8��իN�E�y�?�u��͜��nwr�ʠP���=ɟ�6�[�f���0v��$���b��iE�Ȗ�od��Ђ���bM͌�$Ƨ��O�M2�����A.Z�V�v��q�=?e� �%Ǫ;�/�0�,(�kd��p�=1K�3�^p�(��	r�y�Z_c]�s3���v+�Om��hڄR���eLǓ6��e0�ܯ0/3��V��/N�����(.�K��y���m�}/}�ި��u�ZW����e��c̓O�n}��L�Ҡ��l�W}	,��[~�KL�ukȲ�}�� <�]STm'�t�@��h�%�8�oM�����Mb�~9?����-W�wr]A˥�D	���m�&`���4h�HJ@����ܴ��tz���Iamĝ-�I(t������o��%�_��dI���'��?����΅��3�z���Kk�����P�q�.,(��XR ���p�/��L�	�=Ġ��~x��ih1����4�jA���A�cZ�t��skB,���Bj�\7���T�e��q� iz�lZ(]��>e����7V}'0�',��M�hj�!��Ή,c$R�+1֍��o G�r/�US�Ҝ�N���©adv���W���{����d[�Њ�9r��h�3<qQ������7�ɮ���!ܒٻ\=Sd\~]�x�ÿ�8�x��@Gʊ!��6�c�YҮ?��Lj.�Ҟ�N��U�ђf�c����~k,~���bۘ@p2�u�#v�k���̸P�i3F���u��j{j���big�r#K�n$�2X��uSBi����׾`������K���WO����h{�
T!{#�ս����|������3 �I�I�dpp?�9'�>}����r��Q�%|�s�`nV@� �t���y,�38�2K#�A�k�(]/;�.s�������kb�N�5*��cnX�hrh߀e���UV�\�A�HpS�Sw�o����'���_�~U��g��7�5���d�%�� p�ò)�ZYH#���p��@<8�$@��aL~�&�;�����z|N��^L��k�(!3)�%d|��+0Q� ��F��O��n���t��P��n�-7Ц�E�@C˟,#E�9�GMY}7O�_< q��&�F�ܾ���
���@����`����Vx�ͪ�6{���.Hs	A-����I������1-���"�o�V��g�FG�%ڰ1|l �e@�R��4�Z(X���m�h0=	Ok��[kd�oW���čG�xQF�i�x]^xX��g?��������>`����?��U;Z�bq^�֞{u#�Ws�	5Ab��)�UH�d̲"�FCA�%&�{K���FW��\& k]1���&�b/��g�a8�@���*�!������p���͞/C��Ͳ���M[+ T���ՀG��(}"�Mԡ^ ������:Bb�
���\"������d���Y�����ֈ�M�����������
;�j�4`4���2�9O6��B���Y�$��C�1Oe@@�WQ�3��}b��1Y�ʤq��&�c읤a��r�Q�� �sB) �"�a�2Nk͑����BU��c���rY�������h��ЅD���?=:�.Y�]�t���;�0;a�l�>�D���]}�b|��d�r��őC���j�������Z����G�JSV �����(\S� �t���AMqN����<|�s�M�I�>�W���-�nP4����C� TT<[��U�JI�Th0[��"@�`�{-|�����3? ����xb{�Q��[�g����b�����1��r�G��8M�P�0LV��b��h)�mb��L�ÍW�9��4y���0��.�PN�d���r�đۍ��R~��Mf!�n�o)���"��ؚ�����p�`�sb��`~��Q�W���J�5�[n�z���}��t�j��f@�/���O�e�*t��U�a?��k�:3��e��3S�w.���^�jR�����J��+X���`}�����b����zX��܎�!���ʇ�Óyہұ���i�2����5��Jb���؜L�������r���+�����Et�drĊ;TC���/n\��W���pO/���?2�g�i�����4�0�8"�(�.��X;��y�@�M�����-��� �u�h?F��?zr9�:�5!��'��)�c�-l��B��wV���-l3D[s�d�(#&�>
���U�:	�－�+xx��!
e~D�C��i��� S�G�5	�hpE�g�yh�Gj��_��*�
z�2l:u�`����˞���U�#O�nKT��"Dk�nXU:��s-�C��u?fz�p=r��B���~
�sC�4�	��a�S��Щ��i��v/_@� %���:{E��8@���C��߸��l]C>�" �m2-������M���Z4��
�*6�� .f�D��:.N(�`�����滅�Hc�5_Xll��s�g�����,�gR7g�`���*4�(ҋ"��%
^��τ�ֵܟ�1� %��g�oyot�ú1ڥ��詫���u����Z&��4BMn!ej=�7�Nx�~�DbE�Y3l+]pz���m)���B��ՠ(d������d&/��m���&�����,��Y� ڶkgy�}�,u��t��y�g��>�AҐ.4�E��b׌='�쐼FGgz�w�������Z�b�=��u�e���jh��>P�z�&��z?P�\d$H����"i�B��N��U>��3�K��Ê?N�?W�6�Pَ�%:w���7,!���`���C�[�S%m%g��;�����K4�*�3�z���_Fr�+�0�殎�ޭ���c�[$X���O߇HE<��5'���c��](�.���;>��󥺱��2.q9>�/g��M�D42A���^��/���ѿ��&�wCڸ*^��OG������
�>ltB��%�ٳō���#����f�����A�;���e�)N*=��,�N�엣ȑߵ0/fz@6���T����{�U����l<�Y����N��y+C�7�~>p�b�sQ��?S���QuIO�X�#LI=�KޙlJ���d������y�J�a�`�ɾ�M�?�j9z}¨�
<�聻���/h^+�g�|0�)є��
cUd�(3�	u��^%�17T=����?P/D����K�QN�{������`=�)�\
���iy��7#�·��.;������m'w�8��߀5��;��bf%�N;�0|0xơCZg	��w*#��l�t�ķ�Nq]hyKF�
`_����Ɍx��L^�+�z��/�7n�̭ɚ �/���yW�t?���7 ����'�X#n�lϑ:̹W�����LBڊ'�F,��Ƶ�G���1�z�N�C};}��p��^���a4}�h�(*�YZ���2fq��n��6 �rY���`?7�C�Ǥ�Qҽ���ָ�g���zH��R#�>}3���V(����V� X�K��ob*z���n晠��A�?���Lp�"X�ͼQ�Ύ�S(vǢ)��ӄ�s��y�e�{f�ߛ6,�Xv�I/��)V��4�,>�ʋXV��!_Tq��Rȸ���Ov��f9�I���ַ�Ở N:Z��L��(;K�"Q�e�A�M*@Y�E��t"$�X�	BB_������]���	�K'�h D�/r(���@�m��ˈ��,����xv�4w|+���f���l!/ih���tI��%p��s��i�W���l���u�D���s(AN�����,ĹzK��Fޠ�q� 5�Ǟ@�{dX�,��C��w�t\����6�s� �O,�K]��`�����Ӗ$iM�#E�+g0��q��?��~�tx�����'M� X]�o��%������i?��lž�9XTGR�Q��GE��?.���x�{�֤a_&�=��~suI�/��-hb=�+�\#�הN��*TpFgR���@,�����cݒ-�.�$����Tv��L������ �lD5�W8b��O���),� ��xl��/�	x�����
s_�vڑ m����3Ü��J
BL\�K ����ˠ�{m퐼J+zcj�-n� 0^sAI��E5'�P�~vOF&��й�X�&��V}�P�,�d�wjfk8��;��R!��-|�����c$��(��P��%�,�B�Cm5��t����gFH�a�u&�{z�`; 4-��b�gQ�{%��o�d9���������N�l+�@�.�#�:mb�c�^� r��h�V@_�`_�i��pg*"-� �X^�Զ�&�O���r�4t��$�,euP,ȩ�έ��-�S�$�>{�n�ڷ�)FSS��|�D��+����N� �G�F)��?��F�Ŕ�ۥ��t�q�zy9�U�;d�4g|��B�f�ä��heA��I�6��	�nP�����2ɬ_5u�,׉SB�LO�N�h��oL��X\K��+�Do�k�:�B���N���l"$hD2>�[�St���*yͬF;��C�#&�~j/��Ѧ/v�R����迥��o\:��t�����|�����0�����q�R ��-G��$�n��96�� q!�����l���
��Ў=R=.��rd���"\�n��*H���C��������E)]���l�����"�����A �kdB�xƂ�1@�.,?50��]U�h���^�eg!],fB�l�TXϹmf�.�κJ�}5��C&�j?,����xME0}�0R��_���%�}y�w���9������1,�x����d)�1���s7����Y�^i�D��Dt]j����ޯ	���p9�m>	N�ɇ�G��,�&F���[~�O��J9��Q��{w����� �!!r_j�I�E���x���xFa�A�⎮ٽ.��5�f���T_�;,��=�������*3����S��0���-�K/L�{P�����<�5�cpT�Aa�%�]��C(�7�����nE��(��O��R��G�Ɩ2���:��b�,��  Տ��UJW�v	�����Vx�a��٦�߃<1��I�ڋ���7�=���w���2�]�JE�<Fl�;���|3��x��2nFz�������Ua�Y�&�ڠ{܉Ǧs��vM��\i��t�Jh�!��|4Inz�� .�AWC��z�p��h7e>hy�f³��8�\6�o�m&C{ ��}�Q�]��h	���>]R�<z�%�uVz9�h��ܨUK�Fn� �#��4-=�"[�r��N$�Sw�?8�ONw0C��ʉ���Wn��<?��k����y�r���p�z�Q�4%s��sߨ^�AtK�j�k���/��u���̺��W2�T�Y��ѿ��,�%��,�Q;�)��jEu(�ʴ`����'K\{���7k8e���9�������*U?aAj0FW�|o��j8��K6<����pA*��t$>�J-T��f^�O��*�XbD�z�I~	�r}���^�{��U��W��gW}�MʟQ�!к�Q>�)���A$�����{8�_�TM7�8=�M�/y�����[�W��$�N��U�]Ȋ�N��ЪT�º�B��n��Bڥ�=t*d���Ŏ�e-a[��~<����Ճ���{���f���^&��=��͖�8��P%)�w=LCI�;�~��-]Q�o;��T���g�â��Qǃ�T\ⷲ�'������LuB#r*js+� =���\ڸ�����[%��A�"c�3�5��! ��E�=QC1�g�1�5��anx�'Y��I�<=ޣ:9�8���U1|I��!�Ƥ�绸7���C���&}�9X}�C(�h{�L&;��Vy��ŀ���hn_Bb���B;E~ ��&�2��������@��D$:�B}��0A�w��3:L9h�W嶓9>��l�
=�V�=L�E(O����6�%�(0En~��R>�a�s���Mѿ��6B/�O�n�F�0��7��v-֥�K��1��ceN��6�Nw��b�Ox�Ƈ-Zq/�m��C��
ZȽ�@��id=70�	DN�mX���E����E���>�/׀ kY82K-ͧO���`_�~�!�ە5�U4�^?��T�JQ��89�w�O���=�]�d�Zo��/77�ZPQ�נ`����Td�R��x�c�#zC�H'�&�Mߏ.�M�G�w�������m��p����=^B���U�
K�[U��ѱ��-�T��q��"ã
�}�u�qu1���?�?e�`��6Ɇ$B�5��{����Sq���sz�����0��F9jQQD��k�{�Qs`��Xu�烊�qF׵�ƟIg�`"VDhr��v�5�h�eO�|��G:0)�zM�wj�Dບ�q���|10�%*��"�RG��8n�Th`G�z�t�x�����t��/&��o�(e�e�ܽ��R�"��%L!���*�DsՃ{^D�Y� ����/�pl���kZ@�`=�&RrkGhY����w��BVB���f� ��pI�9�5��BR�>ZO$��1��*�1��Dg?��w�C�x���o0 �@o[�ez�~�\��B��4�G�-|[U	}���W�jFR���b���0��EM%\E,,w�
,�E^���(��x�3�N����q��b�g5*�tt��w��e���
��v�[�@�˖�eC��j��t�|ݾ��������0��w�!C���~p�\D�U����߰��?-�%�RI�����"��="�]�]-�'e���	C,j1RE�{�aQ]��_��aq�p�G�`�t�;#��Ic;FrT]r�#��P���Z�&�;��8�mZu)Λ^or.���N�YG�es�.O�I�<��I�����"�`7i1�v��UCF�c�������t�)���p����7%�M$�2��$ˈ�C��x6m��L`�*O��&&f�1����2�2��^��۸�֓VA�HLԕ�\�T)n:�^vXe�-&�>>���lE�NJOD�"�)5�dE3}���#�+�L��,s~$~fl��5w��jwv�� \
8]�؝���O��8@���|�u�Z���$�z��E^yj��F&��sx����)xy#�g�@eC'Pl?gZ�f���G�� :'��~���QDM�U��Q���G�7��n�gE2f��K��PJ�ͽ�<!��(n�H�p��&���j���1��n�%Ԕ�X��>e�L�lY�vBq3�=��P:������~d�M+��o*I�%���� �9Xf w(ﭲ�x(��!��)
�|�m8��?��4���i�.�\N��i(*�G0�)��g�#pN4�Xn�xq�r�;�c����>o.��O��קt�ߊ{��S8,�7_�E���"=�} �r2r
��N�I ��'�
z�b�Y��} �b�}��몉�4�=�r5��k��J̤��)�-l��չ���]h6ڴ�)���͓��W"�����x�,{KY����������B�L��N����?�z�*.Րi�����b�6��Ԉ�bSD�v�?X	ј����G��R�!����dT��Xe�ȇ��z��G-��a]0d�$ Agߗ���������)[v���-��+ҥa�f�J���0{����Rd�qFkŽ�1�B�j�1�p����k�+���\ڌ��d
^�.����Hd�-�������s��q��0��N|f��J��5_�ii�=P�C(a��.�=!��թ�cZ�Q������W���J��t�mR�0�uƓ�
��i[��p�K��[qZ�e�=z��s�SH{ԥ�.w�q�O�jQ��$������Ԩ[=\��nN��ZO���1��pO�L	�&M�~3�Ə�=�V���v���1��*�g�J�_:���j*=�3�����"����2$ �J�c W�3��Y�Ή~6�(\6������:m�$����L#C<�����'��;��äɖ*�����kL�^&4��n�������ߨh)K��7!�(D�N�p���`�����H�_�(&jZ4�t71`��f�����0zF� ����iN4j��A5�Eܴٮ˻v"�����()hS�%�e�a��9M�m\VwJ̌�v�2�Ge�/ײk1���S@��a2r��ӿL�H���!�ڳ�b��!0���э�����$t�Ӹ=J?'�/�L�􊘮��ӈNC�����,v!Ź������O���_�P�:9���{į��,�H���5��S�$����<���	E��	גL�˔o;���4�c����K��&ȌNQ�����跢�D��
���++\	�U��:{<Z�-�z�7�t.���S9�ze�HtC�s�΢ʊY�V�,��EM��!�J�˲Oc�#I¾a�3�7��Ɉ�wek��Zc�)c�4_�v�� �ɩƗ�av���7X;S�ja��'F�:�1���57W�;�IK��)1p��gcѡ�V]��u�r2���9]�Ƒ�q����#9-��Ӹ���Os�6~�Νz
�~�2�"���[w��*<$��p��Z�NC�'�`�Xn7��q
ָ͆�>�_q$n��p�'dW.sVM?�$��PK��s�Д�	�c^�J��3�/���p�vi��?�_<�섌�E�R�<4p?6 ����B�ؒy7���	�&�Nh�+sr&�Xm�N0-���'�N���C^Mm��Q۫�_�4Θ7w�nLH�4:�>�8�tD���<1��ѩ62͘g*���]���bA>^s&����#-9��,��Vg$h�_c\?3P;#���w�0��[ ,/��f���Z!����	���a��P��+�u4���0��e�J���K0���3X$һ�0k�d��㜞�����s���Ջ�z�rǲF�5��ϧ����g��6�����u��J#������绨~u�VLWU���wxy[���GFq�UY�|�$ޠ	��7�6��� ���B��nJR���`�,�r00:�^��;��{��i$�����4��iD��I�3#����m�l���93p d�{6\`�Ҭ�n�m���"{o@�ѱ���s���W��KK� h ���Z�P?�XԱ�����.�.��!�@1�-{�b:�͎U+�a�;~
�md�@/1?7������a �u��$4�S�!&V����]��a\g���D��im�u��8��*��[i�ne�dD�XK��i~��Pe�O����$٪�)�W�]�gD��a�	�2ZIQ3��h~SY����$<��:�a2||C����A��f0z�Q�W���[��@r�M��r�}�ˌ˃�S׆rPy~�� ��?�_�'�!���حd��<�h~6�:z�Ws�)X���Jq��$��A�ág��v�fNH9����t\~�ɳ��Z�KQ\�%�������@�u�l"�O��.N9u
�v�}�-�{��f�Q��WY0����z�9��>k}��T��
TCc<p���>�}�o��~���Pq�@��N~��T�����՛�\ep��湑q�p�z8ʹ�ŗ\�=TՐԕ������؃_�:�ؐ�i�6��^H�|IA��|&�E#ƨ(Y�Òx	/�Ɯ}o�����뱇l��/-�р���q�N߈�.
�pc������_����ʲ]�i�j��Q-�9��"��M���	"����}��B��w,Т���J ������y�dt�N��5�Q~���P|Ď^W�����e���E�s�����)��j6�KvS��M�%�z7r�0�: -�9v��<I B�fa�����	���Hh~2�~�'V�.M)���21Ɩ��/�&�'R1�h5���c^���Vɹ�%3Y[�͡t$j��Ir��mt9�נ�w&9�RW�Q��9��l��뤱L��|A؄�+I�� �
����@�t��wO9E!����-��{�_>s=J?{��@�ef�(���rw>)����F�d��'*��Byћ��N �i]���uO�;�����+���R'Ƶ�(3�Gs<��H�f��S����~��%����Cٴ�}<��Å��C����6ў�o:	���_�!����(�s<alD���6َ���$��<]���R�%`G)�-��a�4�,������$���'�k�QDg������Z�t��������S�+���=� �����'���H���2,��ܧR�h�-.�.�\�w�K�S��@�^e�Y�~�F��ӞY_E��rp��ӽ=j?HC:��צ������Q��돋=lKj��c�����ՈŻ��_�`k�tu�cV�3>��\�ն�}���-���j+�.������Pӝ �Hn(��]O��� �P6���7��.+eCC���!��h�8em�
��D���c�FxC�cF�gR��e1Se�Z@��S��G��$]Q¤����|ʲ~u��AGB�^̹�u���ىu�Ҩ�<r�l���p*#y�ӱ�L�(�:�L����Av&�*�1yG�:c�A��r߱���x�75y��	E� ��'���_���A��@,~*�÷r��*�Nh��!A���@Ttc���g賟�>�ȸl
�J�z��Ge�4"�(��
���Z ~��� ΁pE�����U�]�MYК��\W�v�N>�o}���K��U=50�H>���*L�7[Q~��Oț���(�G�i%��S �0��((�b���F�#���%���j;�u��gݿg����$5��EBM��V�tQh�4��h�I�*?f�'�ֵ�Y;F�f����|WY��	F��s�$��
�%�V���ڥ�|+b��s1��X.q�pB�1-0f2J�#�R��3Շ6�~?%Lt
�?`�jJ锂CLsV��D	_Ȯs�_�C�en�HL�l�P�.1�DL�d��J��m0��X�)�/1�CВL���������+Ck#A՝�%��ݭ�
I���_���k]V+�lBo W w�F�����LHP6w �����b����#Tu��<��Ӝ9Ҵ5���.�UR�ͣS@cx�Q����vP�)zvp��*Q�Uh�~��\�h�Z?��%��6�[�d4�E!�����_�����Tk��"͕k&����ZY��MeB0������d�P�%����uX�R�����"�O����u�Ǎ�]]�(3S6~\���7�p�v�g�PV6 g���4��i ��Ν<�����=,�1� �*�i���&N�J�B�f��:߀�Բ^>�DV2�y�����Ɍ�\�T����O������Q�r�s)5��/��ǔ�\�燅]��p�Fe����.7T	7�M�˂��l�-PB`���ސT����o��0I�����%S���Q�)
!㧙�2�Ḵ�NBZ��YP+������M-kؾ����@]oqu�"���=·�� �1���s:�&�Ñ
!F:���/,6�NnH���!~�Y�%o�l3�9k�~���ZY�CH�⻕!�J��y�&�3�
���Rx�v ���$FH��f4\dejW����}�V�U�ƀ���ev����s�
�xT��RFRF�)%�>��=���AZ*5Pt��N��YI^݅��S���!�Q���ȻļaE���c�i=&�Q�]��������"��i
�L�.�A7B�r��N0�����{�����QRـބk��K��+�^g�P���D��Ŋ���Vb�����M�KrдhqX�M12�6xZ*vs�U �������Ͽ�~z&��%��Ao�ٽ
���C:���ѹ��97ˆK�Uԫ@o
S4]߶0���]�L�W%{~�}=f����o��=�N�5���E����]��o��v�)�]������+��	��뇔1�R?/)����o
���
��-(���p�齬%+�ӣ�WC'C�g3��j�Ɔb�=-������z���h�r�ǆ��/��P��ޙ@D4g�R`����H�h-T~�95�}����*"a��OS�Or��A`�^y��9e��;줃�eB�4�x�ЏH{�����1�����#���
�o���)�^eӾ}��wn����N�τ\<���<C��t?ťW�Wsw��j�3�`��Sq�����l�b��G�&=�+��w�~�=r�JB}�3��T%�9z��o�Il�l/gԍ�������4���ŭf�j�r��]2*�7��ej��;���c����:�مS}F2��nP?$o ��N4H�C��wS?\G��X��$T���39��g��#�h�dĝ�}����k"�7�~u�a�B⠭�U�`@NژS>z3`��(�:�%KI�?D ���$2d�;ꥨ_?��=�$�Vhp�ܘ�XaHs90����E�+J·P�9koL3���:x�"��*�m�B����Q�o<Z���q'�7�:Ѐ����d�ke�C�&q�b/��n�R-�v�/@�2t5Xf��/�p%�)�P���8Փ�Iq�Ȟ����eޗ{�R��W��xGV+��QA9� �=�E�
Y�"��:Gtc~��U7�(j>,�zC���
piF����R�� �>=}o�։4��ď��}%�%�� .)2��7wI�翮�����̋�dن.��]��a)�Mp��קk�\�}Ȑ6hO0{�����kE9������v50��I��ᧆW+T��R�m�U=$^ɲL��~�,���(d��'OsZ�ݥ�~���� _���~3hh�o���B6���hJ�O�Ro�js�D�B���8��T��n���~h�^$\�n���)���!2�K����]A�����f�	��5̒����;��!������F����Isd�B��L{2F��BY�}\���_q?�-|���|$�AL�L�ix�W�� ���5�#68��������aQ��N�ze:Sl�H�d�Sb�qZR3u4!�#��	�_��;��V�CR�"_���J4,��uܥ4$���QF����f�֔���k���4�7(�Gx14:q\�E>θ/�6\����]�Nd%��1^VM�(td`v��t!Cb&�M�����-���]k���rR���c��n��z����k[y�pY:�,|X���3���O��e��O#lg4���t�<��uP�k���"�H�$�����L�¨4���F�bRp��}�Y��o���w�]�1��@�����*�;6�$S)��u&�J��I11��`�>3׾��w���p,�3^L׈�,��b�v��'=8��:1��?g��k�j7���оs����l�2�ӊ�Ֆֺ�V�Р�g��kh��O�_�����1z۹��-��4�~�E.�Z��fM�B���1����Fu���vy�ɝ��
���LR�*�v�ѽ� �#@Яk�wɉDe(gD������{����O�6D��'/�G�#�q�e��g	����Y�T34ɿ\3=����7Y5��a I݆6{�(��A�xb&��/�Ѓ���)x~��6�J	��������du�ԩ�?����x5�`u�
��mL�K������ҹJ�(�4�Ů)�j�{��kS���Ь�`��'�[{&�����h͹?��4�%�x98�~`�t!I����2��e�6L+�f�]sW��lO�� >��W?�[Ő+}u�l2a�Z��,��b+*�!��j�̒+HZ�_{��۩rBx��؁��f�`X��'55AB5SL+�ܐ���]\�c�ϴҹ����5 )��RlԛO��ĻK��;'ܵ���T��!W�B��Þ�ȣH.m�%��w̢m�E�Fy'�9�w����0�L�v����)�B<�_�R�,��8lk����h����j��뇖z���g��X�/��k,	�'m��Sk�l@�UE�@>�U�~��*~�������\tq�9v�W�{�n�q�g�+�.���dO薽�{hOPo�_�~0��3|]s��P��w%�KΊb��9A������3��D�GϺ�Y����o���Eg�i��ӯ�z�`� ,�w�~����g�F���S�u��w�`�=�P�Dv���]~�uU]29���������T-�k �'*�K6T,j�y ����b����0`fSe��57k��{���4!�hS#u����Vs&�,�JW�V-�h=���g�����N�v�L��ڳ�9�rtũ� �X`�I,.~�m�純�a� lb����nP&��<���ٻ�U̷A���9(����ӗ��r������P,�;n�����+�IT/�hdY/\`_����@[���:�螰hkۚ$7)�2�qߍ��#��RIG�拢�T��]��tn�3��L�T*s7�ڨQ�P#ܸ�ܡ�ħ���:����� �>����ʆ0�!�xR����S���ݾ���dP7�Fr�4��br�Y&*L�ՖK�ۭ>F �'�G�LOӞ�o�1�N���s�3�������,�[�^ѩķ�7=S�T�~VOt"�u`5�$U��T���IM�(JyK���De3].���(x)��� �=�#^ԒH�;��Kp[�i�-�?�:c_�ʏ�����P� �cS:���Y90r��GP��i3� /r��&����1Љ��qL?�.Դ��mp�S'V�b�O>�"����E�"�}��67֗v�oq�?ѡr��q�������=�;֨�H&}�S�QԷ͝bEc��v����^�AȆo��?�*A���� �q��'i��7�Y�t�������F��-j�dh09 �e6#��!������d�7�|�j��}z�	R�b&n�����Sh������5&���b�����a�q��u��f��3/ �m?�R�т
��J�%�r�́���w�%Z���> ����pvu���]�1z�	"{�*~z'rΨus;YZ���T-�C�	Fn]@)�vD�"��JԂRچ�ݝ쮔�б���Y�����L�&���ٰ6��H�K�Ǚ�Z��+�����������J�$�2�2�,��F���4�*��t�8��G��I��Gtl�G�N��Wb��R�K�4�B}G4!�쒣�S#�_WJ �{�9�_��
�t����+%���`�l�|'���X ��B���b�oK5
���y~�3��n*���G<�����՛+1z=�DY� ���."����ϭR���g�������\����游��p����QǱ��s�f�a_-��ؑ!m�����g��u���hz��O�a;�&����u&�9bo���^��{>ຌ��N������0��� �S��b)����i!��$�'y;\�R&��;���Ut�K$�������8��,9�|��pK� ��w���w4޹��I�S�R���J<h&�	���Q�C�9�w�~��LC1''�j��(�"��bW�	��cz�5?���O�:����:��l����J՞C���[y��o�P�$��-�@�c<ģ�7�G1Ԙ_��0���cF|�*�;�$�2��tܔ;�˾��g��;'�ZSԕ��k��3�>�Iѐ+4l|({�w�!Ŭj�('zf��ym#�ʉ~<�7��A��(��@�I@���Y�#��`T]~.�D��JŕA{1�:�J|D��t�}q�f�s�����wS��|L��]��ai{$��s�M�\�EXX�?��ЄY�M�m����l�z�U[��T�ԗ�3Gv��?�@ ��k��;~�/U�hb��}���Z�SY�sE�TP~�\ �jɬ����R���w^S����e_�d�I ��c����̹���_ж7q4����
`���=^��0hAdf�fxч�s���tr��@�D|��b�Ǆ�o%-I5�j̬��"<�m�t���J���>�>�~BUa��G�"��3M�П-o��Qg�w�WkS
� k�z�[g��?sm��!��b��-��^�qCG��N�<�!izQ�wY"�:� 5`�����W$n�I����z���0jFA���X X�b�W%y��rx_)cQ\Vd�m�7R��"O�s&��Q�aK�D{�-~Fi���<�3�đĲ:yǞ]��GWNs�ȁ�P��#O�a�CY��4��<�[��c�;K�����M��R`��*L>�j�O���d��cnGUy�ˮ7���rH��D����h�
����U�a��O���?|��A��M������{��N�T�0[�w���|:ͥ�ZQPM4Uvd⣺�c�P�y�,���� n��(�U��/K�ك���i�|����v֊V�F�gc9�C�p/�-3p�^!>/�-�����C�C�oT)�h@N��5��"3N�&��l(��czI �ؠ��(�Ch��˝?u����Z8�Si:�T���>\���ML�'x��eۦXܙ3o����,.���KCa`B��|�B��4����P���a����lȳ����x�X/ �0Y���OL6|w�������e66:�ү�	 z����񝍝
�v�]��U�8��Yq�$��m)��"dc�ɍ�7���/����e�4ת�h5µ)�t�t�Z7i����i��/5��e5�Ϣ�7�n+Pl�?��2�М$,�>A����H6���aaq��� Qg�V��hh�~ EA��Nj(��R�7�T�vUg��B`HK���c&���'R�ED�c���՚��𶓸v]=l<���N"й��*�T;~�o
=�3R��� �� �O��|��Dvt&���=�X�bc���_/�&u5��g�ez�����e��!	Tꋊ�'��;�/��a�BS&_g֕��,-�]1'�͌j���:A��p�MW��ZX�iγ��c,��kE���7�k �(?�fD��+[�F�V.v�w-]��	F=asǥ��ӦF�C�S��m����#����Eϸn��Rz;�7���1��P#Ϊ�I�Qv��h�ݴ�oYM$��#v���^~�k�쭲$9��u6;`�4������V@W��?��V���������!	(�d|�]t��h��`-*��T������f�p�Ti���D�>�Tb޾�������h�_R��;v�)r�(HɏZ���/�r/J~�gv�x(�q3��n���	���0%0&௑���yU��I��0gD���l�]DBL�b�Qx>ƫ�pP��A���wtPi=<u���LW����t�M���֍*U����%h\�7Cq�!O��d�(����s� ��o�.�F8�RŌR�ַ���!�Ȩ��Jk�gQ��=n�l����N�#ᅭ�A�͵p���}�s6�bn}��~�S5?�BO,+��������-*Hҷr�������0j���E^�Z��4l�ԑ�2��T����՝2����c;hh�ykL�b�9���P#ABX�$�
ik��9�@
��&Ys��*f�:)���Q{� �.{��;�$��m��R1��̓�3�Ɲ�5�JD�:<n_��h[�0���2%5���-��޽��UY0�;~ V�Ȟ����L����X��h�^�]�Nj��4��_L#R�6�g�S*��03Kf���!���o$s��U�3�3���L]�^\U���=�X'NZ�v�
��`��5��`΋PO"Y�=8�^�d�(���i:�<t=�
0Z!g[O�Ys%M��w��\�R�
���3�]��k��<�{߯�hc�{�d��ջ���T�tN^���S�L�۪�e�b�PÚO�ĔJ�7�_�
���س�Ym3�t��6NA��cd3{j3A\G�w��&�Wag�
�Hb9�d�mD����$귘��Q���2�
��@�3bi���`����Sz^̺fo'd4S���ٔ��ā��Z0�P�f�;s� \$�6@��K�L�Tb.Z�����F��(�˪�*X���O)�<���X�W�@s���S#�!���-�D#�t������a���gԞ�t.���t�]��l�a������}�Y���W���rH�18t:�xa�H���zd:l!�Pta {���mT�y�6�^�Ͷt��.��q��E鳗d(�Vو�tje�J�Y/tH�0�Ja���=�ƣ	�����{���R"��b��z�¥08��_�O+�ϪG5AiYL/�|�vTݻ#�HW����e	��/���)�lP�c8�� ��_���'K/��h����L�>	�6�D�	���]� ,�95�Z��F+A't&����caGU�c
�����&l��b��fq��s�wG���4���S�H5~K�Z�H��<�D跕��a0z���l�j"Kԓ�}���m�/S��˄��Fۦ��Ul}#� ��!C�Î�p�׿����#�%u����wY�}�6_`� �݆q�Gm$A�~�V�
aE���ڥ�
�M}D|��c|cT!�IeTy#�@+���}��\F+�Sf�7�/�O��P �!d������(��\�9��jӹ��a�fZ����5�YD��Gܽ���P�B-9�<X�&kB6�T�O�
e�[$\�õ���d�D�D�^�`�k:#�)����x�-D8��ϩa�I�d���q�f��_L�ϥ��B�"s�����.��82�Ę�v�M&�6T�c�l�!�} T��b'y=���0U�S��i�h�<^4���郺/��ƥbN�m6��~, ��A��0L�LԉG}�d��I���K͌1U?��W�������*=��[�S��@(�P��3��=����z.9�-��$�$~e��xl+��>k�L�G�=�b��q�.Ŋ�Y;Ap%��|���1���re*_^0�*��B	��R�
���)��ڪ�Ңae��P�9C�뚺���VC�g��N$v,|�>�rݭ�}�@6�Sm�f�s���7���H[��:O�8- �!|�1i��8��\Xor1N���
��-/�_��5����EJ����<j>�����1w�ld� ���,�������_/����A,��O���3� �hx�}�gn�����Rh��2��)p�LT� (�be�+a_\�ȫp4w�ZMEk�m��v}��� �*�!�O:�A!�UԤ1��cN:�c����ퟔ6 \E>��q_"�a��I N9�T#	����E'�a�_��a�h��j�����[;�g#9�gz��D\��u�U*��](�7K�j���6B.څ��(O"��ȋ�(UMy�92���>XV��,�Ê/q�"�μ�Zuj g��49)k�ZTh�;[�/Q�@/���i�����[��Nc��Dw�Qmӿ��0?k�d	��f}��5nD�:���"uid8�ɿp����u��>L/�֍�����QB��&Ҳ���δy%��1J���NX�Y��ؐf[.�b��#L�l�c���-�6� J�M���T��V������y�T����w=mb��k�Ejz�3�w���V�kO(qr4;��[e�������X��aMKK_Vq;�-�|��)b�H]�9���v�a4J�$o�����iq��+���?�_�)�^!a12��՟]����:�L@���F��<�D����ԾOO�c��_>X�S[��!!(�� �b�Q8?�m������&T T�7we,]���_�䎌L ���g���,�i���8���*��6������oF^�8L7Rv�l�,�ʆ��;cx�@~5�ZP�״�q�o�;��j`�v��A�Qb+��- |E]�au[?������ sՕ�2�����s�2�	m�U�FP��O�����E��K���T���{ag� ��#����骬��;gLd�z�zP�����%��p�*H�'C&�Ϳ}͟T�_< ���$�֩�>k�Ob+<T\���r��%e�6	a����m�Ҕ<xB�;ކ�\�7��hֈ.N�p^�@`�b0Jr>1�Q��]-��g�x.��� lMc^=S�R��ɐ��
8MA���ʄ�����=[H̰�R�p���u�(��GF�J����(U$�[����G�(��ф>>��O�;K���t�l0����K��ȕ~��2��)l0'�%x35Y����O/�����m����#��e�J�C��х'�GU�в�Ȟ�z��o���'f}t^�zu�h���$N�y�R�<�����K�m�o���;(h3O��f�B]�Ɛ�a����h49�=����U��!=8	Y��0\&xop�0GNY��p���5{���J*K�����m�����������W�����`�d�5~�;�2�WJ�o�03�̥ahF�L膞�/&ڒ��/m���j�0���vg1�a��Q�B�����&���!^��>R��%QݳA�`��ψ��<�N l7�|��$?��]��82��-��,�j���=9}�mD�)����Q}���/�n����L��yZ@�kH��ٓ4�aHEu�X}�6p�:��pZ�1�ɴ$�w�<���f�ں྘X�VJΦ@n;o|�L�L3�5d��Z��.wNln��!b�Kks��S�-��-��&���e�(��RQ6A�U@P�UU��<��Q�x.a�R��EPc""���٢2���-ʰ<�Y��ᣪMWv��ҋ!�����Ȣ3�T5�ң�[�u,��/fF��=����=�OY�C&s����I�ʇ�g�}��D9��Td�]���	�qƾ�����36ٍ���s�ӊў�U=?�_��dŇY�)έ�Y�Z������}i����J}��P6�F
<B�^c��l��ݸ���Y_1�sV�dh.@�f���C��p�84h���-�S�T:<v�h���6oQ���XE}Z+�Uz�k�h�?s=�{3ֽ�,$M2d�#�a4��ݚ��'-c��oʍ���o��h�[/�I��f���Y�-������y��rU2���p)-����,'B���Ot��e�ɳ�	�s�Rk�#[řP�寡:[�|O��4� �P�h{��k�`_x���c!��-C��f�-�H��l�}}�C�:R�ַ���=�Q��'��s���>H�r+�Wd-��$�&Ϫ����]�詬Ѝ0#�|u� ߴ��9�כ�^ p��fG1})��GK�����x,�C�A�e$��y24H7 �[��'����U��7!�k�(��vA,h�z���Sp���C��P��
����t�9@|�SLc+I��Z��v��'���E����f��_�Us`�S;ј�
�����G�q)#���F՗�� �q3,T�9�5���h���,�b���i��y�AA!rZS��M�ڀ�Z��;���L�-���<��`"�]g��~a���R{bE�:���T��W{"%�)�~a�*-����{�\I�~��~b���Ċp�{yc�d�Ewb����!��f�e��ؒ��f�@ݒ��>:A�xQ���?x�C�E5�����a��o�``�S����!}��33at��({#�;i�i�t���|%���d��.�}p�dޮ=��N��G
����UdW�_Ǯ�|��*�h}/��D�wϯ��˝��2��l���9`�+�=��܋��ɁȿQ��]��2X��§���i�����6��^��xw��+�[���Ĳ*x�� �I��d,��`O���{:lT�n�=�/����9�s�T�����'N���΂�J>q�ܑ���y�W ��C�K3���������e���m�n�\�oI n�r��'��q�{�x�:T��<�%;�zSتGZ��J�%rS��.��F6֋\y��\�?*`X�0K��!j����x�ѹgB�HS�����`-���r@2N�.i�ĪK��
��eت�@*=&���ȩ���E>���]]�XpO6�P��ݵ����X�a�ߏ��)��v%��eꓐ��E����q�t�^�.����W�4��ڵ7���
��9�0y���g�U#�4��W�X�2J���`X�fl���r�P��`9Ty�D��g�D�!	=# ��	��/���t���W��x�7@��L�wTs���|D��F����T��8hX߫���2� 0? *���U�}0�����P���Q��gPV_Ibq��0�j�"mٓly��v����zV��)!ٮ84j�ɓ��q�s���_0�tz����0�DF�0l�»�B�U"����%$�/T��#�t/"��v�_����~�� �w�/���CB����M_o���< �<[g�� ��Lt�~_~�G�u��W��ˆi^jIg%��߯x����B���E��J����4����Gi��2���)͸�4�=C1B�#�_���d�4T�8L�i`�B37��*I�N��E���
��\eǬ��C�p��$W�4×%4VL<c0��e� �I��ˮ��G�j��:M�W(F������M\ELDĕ�eH���83�&��z�v�ɉʰG�������=W�4x����#��4���(��w�?[̄�r��w!� �Y1F'��@ZӞO8�����x������l��C "<E|��l��?5�,����b���8/$㌇~��H�d(8�:��'��eY�r!%T��,�Φ�+�>��������`1�b��8���G��l�^�(���~cp��?K���\����)0�BaO�h=j�}���C�|V��ߊ)�{�ȴ�T�́�:l�0F���l32�W�P�S}������1�����*��Y���������C�&���W��Js�wW�y�����;R�D�����K���_V΁���߷���`�w���/'"F��i9���� �YRc �AK �G�溽��s�D��w�U$�s��&�_���dm؉3�G޾�+��\Q7��zJ!@	��Cm���v�E�[��*:&�d��
`�N*��}�;���1WQ��aN�$��xqi%*��Ēʧ����g{�Ŝ��A����D��RS�^<Mw�F���l��$k�C֭}R�ͬ�,�qR��0�>Q?����&Y�	��|������.�IDoA؜򆍢�)u�A'�c�e��i��qi�������'k�w;�#���+�7���d��5�.D'�Xrhm_�˄,T��lb��6hO��Ìh�r�$���(e!g��Y��%���Hր�;N̔�hϤX������B���#!H"?F~�a*D�<�V`~2�YC�Y12T�jE0=;��	3�Y�T�f�W�n2��Q �֜§p�� 	K������<m�7�#"
M���v��)�!)�}"?��'V9f�Э�Go�ʸl�G
W���=�.W���"�T):O-nH{�IwT=���go�T���d�rF���#��)�\��%�ޖr(ŕG�&�<@ɱ����Ɋ��ޖ����ߌ�e�b*%K�mK���[���YW�*)���ߑA���Ѝ�u������߯��wտ>����/� ��� �d���C��G�o�^��Ǳ��f�-�����i]�r��Mh�6�p��L�����)��ò�D]��M#���ƞ��)����4B*�=���x�,4b1���nAzi��R�ʎn`��;6_d�ߒ��V��Ǔ�&�u�\ʞ��p��nx�����/W6=@T;��Dե���z�p�R[�b�F+c�nO��f��})�?���\�,2�W��.�kX�u��M!�5�r���l��:��֙�<��{e4�j>�<Ul%�t�3�9)K}�0N���c�TN0W��	n��RX���d_L��",���?�����y� �;�KQ�9��?A�@c�#alS-zU4ײ��Cz�')0�"�p�*+i@$�8y��c�xꏬ��T?#��5}綮�7S�'l�.#:,��F��q����YB���Q��M{U:��3�����6��2�Ӂ�]��vj,����&�>vd4��X�������N����Lݸ�?s?ӸRZ��+�䶟������F�2~���h��HqB��R8@�����4�UhЧ3�;0�'���� <3(��ǂ๰
T��)��oUܻ����0��}���J�z*�kS{)�L����ICP�o� <<@���W���3��`d�p�(���� �o<��&lTm��MO����o] Ks�퐖�
�΅�u?��a���Tu��7���Kj�F��B����iNthQ�n^u)��r�h����aUl
��q\��/ +��ix׬Y]@v�X�'95��&s��-��[�(zSp*�U
#�E��e��$"�E������aG:Kޟ�|��)�����uRl�L����%���a��W�~{t^���Ο�������� �&�?=���J��*�Q/����qR����'IkD�2���wܧ�!\A��<��ƅ��B=�o~��-���S��U���
sD�#m�y�K�.m:�Z�a8m�ݩ�*��Y�گy2i-����k�xԡɃ���ElbV�Eɨ�q�.��>��`��oq�1-�В�z
v$�/?n��t�P㛏0y�T;��'�h��$���gMl�1x4n���P����WCgp9��� ��a|�3S��C\~��dJ8yڔ�a�`ι���}\Gݾ9V;�5�c��G�nX�4�����t�,p���ӥ?���9� �!��J@�t>��ԣ���R�!&/}(fA���V������LwU���}(��Q�w�!���"/c
lp�3��=����-�A+��^�h�Q��}O�Ќ�l]�Xj�{�[G>gqV��!���+hy�+���S:�����d��n�䇘h�ʼDj-�Z�}����`�x��i��	������7�8�zH0_R8X��'�2X"��lN��t��B���I�b��Hw�5X�tz�
U�L��FU�wr(�L��*B�;���"r��$���/O������E�.(I��T�o�AKx�ZV���:�ь���,n��F^��9�3:;�!�1��]�������N~� �a��Oʿ^b|��m�H�-ylou=�_���8槗��_~͑�yƘA&��g)���q�Ě�FϒP=��PP�˄�c�8 'L�Z/�m]���Uh��u��Z�������� �_ۗ�t��RO��C�E4)D�?�ԉs��9s��TX��+�gXZJ~���xC4i��n�����|�Hd�-5l>�ƃ��/�ؕ[n���D:Ő�b	U$:ߘ�� v7����+�p��0�y�t���i�t���Js�ǶUX_H�w &X����5pZ*7�Tۂ��h�E!�����]�Av$�n��/2�0"kKv;v蟲�X$dQ�\k>�@��#�g?�W��N���K)�Oh)���:'5<ow�ŻB ��)�XH?Ӵ��|(\[��[��v��#��oXg��>�<�.��Nޱcک� k����,�;�#Tc����ím�F:��&��<�WxӝJ+����M� �
::���sRfSD��<���;�X6K½C��#�<��t(��Ņ�y��P1�|0�]:�x^8��ƠSrE��c�u�mޓ%;���>a�X4;�L�C��z>��F�T��%$��r�jQ�٫y3��C�t@��r��c�|m"�L �\8c��;���ع��W�=*h��2ζ�$d\(̒�h���#u��b,���4$t�ݢ'�&E��	Kvs���>j~{�9�k��r�H���
�C5���E+�����0ێ�p�p�����
�"����Oy��{�~����g]�Y��/�.E���FÐͨ����U����s®4�S�U_�Y:���5~!�h�ǖ�G�守`�٢k�O�_G��5��s2�P�7,�!�����*?�	5�e�8H���z����j��&}�'߲�V[��Xm��B�,`d��]犉��/����
˖�x�&r�$��}�˷-Ԋ��h�q?�%��
M?4X&l���M-fh��h$�D%���l`l)���7��P6�,!�)�Qďx+�1Z�QS�h#-%��"�׊�j�%=d��������G�,��!(�^_};6�"k��`�@E�fê�V�gP�n0�cP���/Q�����U�n�W���l2�fS��.Ì!���~�|�ѵ�",�c{xūɠ&���ID�
��e�T�A/	���+#��B���C��5���Nu^D�9�xu䳡����M3D�ɦB#����mF&�W��N��c;�x<���J���X-zZ?����E�h҆.��Ew(^��9 �f�Fy��u�6�s���#K,TX-��0�U�-0�������8�kb��T�hn���E*���W6y���P0�H��ΘŷZ���h�4�C��DB�s�6R����^�ج�
r:9(��g焎쬄�;L�����ړ��"��t�_q����
��-��NȊ �#;C1��ǋ��:/���C?\�Ov2��;E��~��GY'F��J��"8�ճ��UM&l>em�x����AT,��8;��	Ĭ'j�H�_�ge�� �X�O����Ԧ��N%�U���pӂ�tRd�ɍ5ΐ�Q��Z9s���<���V�۾DZ}md��˄���tд���v`����d��,����{x�S�bǷe��-o�V��>vJa�D��_6���5D�,�_xXw��a���w
�	5�m'}v~����ߞ��PS�=��\4��I`���aҌ�=�O�UH-�IÄ��.e��W��?���>��2�#�y��;���_wl��j6���2��%�,l-
�Z���_�t��۵�ɍϒ6�f�����f��{UU�J��y9i��&T�{D�Jʬk��Ϫ�Sb]��>�.;� ���^Ͷ�hy4��:�aұ^N9|�7漕{�$�e���VkR0|)� 0��w����^�F���7׭a�S��
����;|��^B+j�`� �Н13��.6"%���ސ�|[�(P9�=
i[�|)1��@�eE1lO�$h��>y!S2�N�
���s���o�Zp��ˬ.L��̌j��6_"��1:�+��96#݉�Lp���ׁ�RpA��:���S#����G��`���X~�"O�ş�s�]+	D�c��Uv�!��s
�%�=����0�s�Ĵ�$�U($`�-�(B<%�P��8�H�RmIЙ��5F�I�����&h�������J�+�`�GW<y�|��׾�����<���Z�Q<�gL^��5����IC�he	��G��5��'�o�G��751A�1�qm�-����@RA�q��W����Y�Ft��n��%�����CGqYq�R�ff�ã��v{�o�eP�W�=�L��_��SBC�&�q]D_�%[�c��w*�C�X���\F�]/d�*!����ʦ ����d�6�%���x���0PX��$!$.\ԻN["j㺪:�DR���� t��C.��� �Z� �{oKg�f��`�6���N G@S���"/������Q601�-��˸�2�)�=�U��BZReȑ4�>�8�s�����=.��X�jٜb��(�g�:��b�u�Aѕ��UO122R��[U��ڇ���B9Q%���'�v�AmX�����y	��W�,�eKDzE�q-���6��?[��81�t���EI
3$��j:��M�������#�%*�c�̍��<������mc�������\�l�Lk��s�;��Gb�q����Y()���`�5c/�;d�cm��ۚ�Hf?}��t�(�|$���# R��I�ɘ{����}^���{3��3g�ݑ��D<�j�OI�Y�������Z2�T��2{P�j�吡!ZZjtH�a
:��P�6H�"�0�>)�	�5�i㧻+n�H!���yѡ��5�����P�=���6�uws�f��@��q��H�ŏ�0%Y���N�Խ����m@dq��<u����(}x�

~����ft��+��&t�X S���k��UX̘?�W�a6Q����<���`&��4���.{6� n�L R!>�N�]pՁ"��>��e@͑9�]��n!"����B˖$����!|�T�����9���5�ï�}��|C��97'[Ԕ9�p)��-��@��T�]ۓ�#����c<���Ń@�/k��	��.�y�UlZz�cw����Q.�[eDjln�hB���~;5gm��C�|�\A�K��d�P1*9vA=>+�B�5@��	�f��Kc�j9J6�*YЄ�)|^���&�9�����Q>�ݭy�a��?0�4��Nʎ�P���>O|�cD��ޣdڧQ��)�J��=�f
G���������|�e�a�`�|��Ҍ��ڍ^�d�i��Db���Jo �	�.�
#2��=¸|������V&��,���T}����^��,�@X@}����4��'̳z�*hҽBf���{&�{��}ױ�0� @�X�#�׃�~b��y)�4��K'Y�����԰│{򕴰��pþ#&���҅ey���)������,�V�)�(�$����Zr�N|�8Ļ�:H������7�VrE���~������cD�q	6�hQG�4�,��iG����3�����VΎR�O\�j�+3xa����.��N$%���=Q��ό�WD���\�销V�
F�%��M`0�y\.i��uR��BB:�O�%1y���a2Ă`I-8l{VӋvhv�@���)Ik�3\�M'����?y	n)E�jg8�e vj����zCz���M�L}_ʷ�������]���q��Б�[
F�Xe�[B���izά�9���]k�2����Ȩ��E��D��:�z5�����O�(�U�&'�#Ku�o���X\DSN�hߣMM��������m�k\*h����Kᔌ��h-��ޮn�ps�}1���l��d���?Jgc�e�����Q�l�v�x���{��5ԧ*k�����qR͵��N)��?K`ٱ�{*�D]׋�r*����\.���p��6�B�Ǣ���;z���TM�ݮn&M@`:fv���RJ��7��@��c�r�q�u�LJY����ܡ���;C-���{j89�X�؉��O$l���5�SO�n�@���������6;��,���R�{Q�=m[�q�Éɂ,��t(*T	)u}�&����HW�.]���q	���V?ղ�GPoɃ��<<:��a������**}�s��%�)s�r�XW'4~O�������d�/I��B�T�=J�?� G��R���-Ţ��d�L��⠧��C
��G�uH܆�0�`g�Ao��S�̉�O�K�~?T���ﰹTh�S��:4p��`��޵9��s�,J���)J�u�TE��X�[PR�&�ZϞ��KG=�Q�Ď�{4ƶ��d�d7DI�:���d&f��A
s�.�lƔ	u+���jh��wl���d�`OK��� ���L�~Q��y)����9���+�x��&��&��Ym:Y���s[ s7)z�7D�L*��$��,�Z�����q�^�{�Uצ�i���m�	�y���l�Vf5tPb���<TS)��7�GՕ�q�n�R*�K��A�[X&�'w���j_{Sȭ���:A��D8_�3�1�Rz!�"�6�X�3{�`i"H�)��}Z����&�\�X:r�+�l���&��;���H�	!��u�x��r!��ë5��G~�U��6�K�4=����V��lTK� �V �Z7p� eJe���i%7;�4��e`�NN�}��(��RG �IۓC�9v�y^ T�&^4���l}�z���^
�Ѷ�ZX��E��5�U�"c�HeuE}
����]E��*G�{j5���N�3�te)�N��Y�D�@߇&�Au�o��@AJSU�0�m麣��� 8�iA��� �w�lΈ��4>�9���<�0��ܷki�	�d���Ă��`�Y0��i�,p2ze�jq'K"����<��8Q�����'�}���9>�JR��#UT���v�7G��.n��a�:��)l�ό���\ԓ����QNÑ�Y6�&΅��;�ϣ���t	A;l�~�"�{���:*�ꓻ���J����GX�u}Eq��yx��v	Ӟ�Ӥ��j�<߭�?��
�8)e����]��F�:_������ߏ��:nJ��[�7i��#=��� ��&����X�p�@�|@�0b�ۮv;F��������P��D�L�nPxI�N�8�X ����q�B��s���������U�X�|��#�ɗ�-�Z"r���d�q��e�i�:D�q)<�dt;~����`�
7�ޡ�k�,(I�l���?�Ryaawlˋ����[�����k����N�B����6�Li\���z�U�Ø�7���������4iZ �\w����C�7]9�l>�y*@R9��	`�޼���������
u�tZ8LE,I�2��ߟ2�S3?�}������و�˨��!c$T
I����﮹�o��867�|��)�& ��GA3���_��WQ�w�h�}ڌ:�/}��5/]ߟ�O��Wvk�u�[���>S\�U�ŗD z��w6-��\�7���r\���O|��GTw���� �&��9�)�KmyqH��$�����0��L!:�	&��D��'�;m7���IG�Th �-~S���'6_"*�ծ���i��ћ�������B����f�1�||���u�u�˧�[BU`��;��S��X���/�/��|%8�M��杻]<�
����]I�p˯([�g����_u&Wd���6`:�U�TR=��ׅ�.#OB�o{�x��w����^���G���Je��t=ҏ5�V7���M�Y)
�8���uLb�y��k͸�ԍ�(���z�^��#�V��M�@��9wRH)Q�6߹Bp#k�����o�
��M����r�ߴE��6��*�0��S�1�dh����q|�[⪄�SP"�e�`q�4D�� |�k��b�֘q��B���Nq�EU3ѣ�������=,��������C�`Ƹ�k�J�~�U����|X��tNZ�3�C�:0��1����v�\1`qB��^�H��wD��QU�,���{e�_�����ET�ݐ�q
�,dNf -T���č����S�nV�A�ok�7'�dީ31�v;��w�W��a541��Y"�E"a+��-����>�ވ���K��a�?s�xl^����G<]'y�0�Ǧ�\�5æ����B؃���������H<=z�0h��1�̢<
�>\(/�N�H*�Wp����	�qΑ|z�e�ョ�� >Y�>�S�.�xٌ��(��9=C�L����lH�`���7^�{��A[�Yn���9-���Zp�~��߸<#��n�篲[O�qԹ���F؇���8f�j�8W���yF������Uc�l����j�ϸÀ2�i�çz�� �b�7�Y&9'bp�SŶg���g�U�������e/@�	1�x��f<�������p�8�I}G��V2�� F�=�����_7��|��a�.V�N�_j�I	��|wjS�O1ӀgxEe}�[k0/m�=���6\X 5�ĺ���-�x�o+*8���*n�������y��? R:�i�m*(���F�:�xu�n �����"4{Бv���pP�M�Դ���R��VX�H�nGDR2`(jT7&�s��)�o{�3�E@M�e0o��l���a�P�l�՘�J�X<G%~��^W����p��<!�������'gͱ�:q7����O����x�p���������!�:���m���ɱ�X�N�]�֯��	�5��I���L�Ǜ��a&�v��,��f�k��k�xB,�o��B!���>�| �-��Y���(�lx�A3�X �x�U���<P��hO��y�hcwrG8�h	���Iɏ��������&ƹ�[����h�P�22wA��W?�?ڭw�PH	9�şm��!J��������"�h�K��"��������� �=�.��0�4y|�o~�~	&��+��؇ -�+��0��Lg^�eW�q�(�'lzo�*|��,*z����"k������Ǩ���iM�#3\~Os[�t�|�@p��^!:��0u�Y�}������[AB�0{�0F�E۾pl�ex��Oe�n������'���r8\�{1�_~�!c��5-�DwN"������ĭ��f���p�U��9Ati濷�|p5���N�Ac�k;��L�a/���<#�v����S3�)��s�0M~ U#r����'I3�E-Y��A�$9�����_e�D��z;^���,k�^s��Ŧ��M�t^�>>�]�bê)���M�.���4�pb�m#܈�b��ȴ��\P~��o�|8���P-l�0������{2͑x(e����=s�̊Fi���y�1B���kF�V؟
��m�R6���,�kN%Aꨛk���2%D{nsn��R_[���)}C�{\7֭S^G�x��~��[ѣ�i�tU�8*�<���Q�؅/~!����%��:V� 
�,����U���%����}���Af+�y�
t�QH6�"�&w�����]3����\���S'7�yf���~#���P(�N}]T��\����*�f��"�}��˽̩[ycQ�P\f�X�� yѪ���:ulȄ���%q��3���������i+)ek�o����|�Be����3�Ȯd�JX���W�p�,p}$4"��'u���jy��"Ѱf'�Խ�D1N�j� l4y�r�{z���W�w�:��k94�k֐^uCJ�����\��T��#N@�G��KM3�ہ#TRj y����&�rW#�h���87�?���y�K��'ì�m7b�ton���P�������N��UJ=����[�T{��8NK��T8���P���JG]�_���� &~'�m`^�l�c�i��Y����䡌-�D혺��mY�b��&{���s���T{z ���.�Ms5�aM(Lp)"T-����A����J�TPlOnO���ې�H�ƍJ�U�/�����FD����+��d���0��e�;Y�G�b%Qj�m�EI��G�Տ�=SR�����&�;�>�F���_�Ǭ�A[L@�}���9���`�����H+�&#���E�&iv��f�m�h�M��)@)�4���K|�}H������}��[�������Q�9ۘ������07��oM�!Vi���i��̈́��&��X~�dI�3RvY�<�`�z���T~f�4޿��HP�{ �D@Y�����+��>�ue��
T�h�t{V�U�o�o�8��sѕ��F�S�t�YU��K����-Rr�#��5	6s5}#ws�ry�!%+���}a.����L�/BYo0E#�F�����J�=�����3���cw���79�#[A{_����4�2U�|z@�8��>�������	���o8ҾAݤ*u�ۡ����2G���&�(x����ӹdB��X�K����Gv�` kb`ƺ0����>����\�q�?_�i�P7?yG��"q��X�X94��8��&"��i���^��'�����%�v�^B^��O����<-�m�V����� n���>��i�0qN�����ɇ�\���EaW9|s��q��|���{�4rS咂�V�ऄ��� �E��y�#�g}��e����Q�j��k8�m� F�֠���	����`b���v�Q��$F�X�V~�������fE&����Bm����
'�o��#rB{�NK*w�#�>G�~�	@�rm�N�T���֚���p����1�?����z���RCri�	�6zY�K�]��C��-?���&Σ��lm���N�i��$W�`��X�>y�&^�f뚎KU=

�����Y��T����x�juqRO�ˇj�����y�B�(���fag��jʌ�'k�b���x7ELq8�'~�=Hh��(�,�g�p[�u�(����������P���'kh��z�B�Z���9����V�y9`�d�Bi�*��X�$�ˬ}$5h�N;���~����*�,Aݐ|��"LC�D�N���]�� �����������y�1�y�96�݌b��S a�SN/f�Ez?��z�5�s���3a½��K���HH(u��c���*�l��bY<����=W�q4�ߦ��]���ʫ2�V�b�V��k���pf���oi]m�C���*O�heШPFY�s �f��֚k��÷W3��7��c��_��3��ĪI,��]�W>J6������p�ܤa�6��M3m���PO��4��D=�QRh�>�ni�ª|�I�V��~H�Z=k��<���k�U-{uS���J������$+(�r�1L�i`�t�2�����y �0U.�"��C���Tmv�(��;-�$�N���J^W�Φu55	�E��^�u
�0����ܯ�d�}��b���q�	�������F�� ���(}�ǉ��"���X���jM�p���[��8?�*�]w�&zK��W�A\�>��-f�����Q��k�<��^��V�������D�k�ʐj`֏ǼI]	x"M�@N B�} ����{�
�Ӆ���\�'-�m?ǫؓ�PB��ϙ���L���VX^T@�vx�O��H5���u�&ʏ1�yp+ �b�0p�.�����l�1h�����ΐ�-9;�E�oa�{0� ��IA��"�f3��1;WJ�ݭ[ï�\�b;�:��/~^���v!DZ2�@�B�+�j� ��В�Ru,d�Z�kX�Bc�S�d�0b҅�o�{�H�q؈VͮD�@��9������@���,�K;�w���l8g�V���-�T���y�BFj�x:��[.Dj���K34R}�n�E��ܯ�޲v����:T\q����� e��؏��\�4���uJeC�j����7m��D5�\5�l�Hi���!��q��J��l�l�}g�#����J��!"��t�#ᾡ�eEu� ]�1���e��hܕ�A��E[s��1�-#_�8t-x^W������Lj��. 7��r�& g���jE���%�Nk:ek�i��|�|�!�-)��Jl´��U)��W�t�D~-�o�D���f�G@X��-nVS�B��M3#�Ԃ��:)�L
��u��f�x��\3B�Tx
�o�@;&��	pm�֌yE���г�Xx)�_�k�37�a �U�0v��̿bM�����x{t�^�n����D��ci��@��pZ��ύv8	���K�
�¯C�I1R���i�̰�N�� �#���J��bT��.�b�-�W�"��t�bCr�X&)Hى�T�;�n��s���C�)i�4� w�^a�L�X#Kg�u4H_����c:�K�(�;���0
8Ip�͂9����.�`�yQk�[�AS�K����qN��-B�>a<@E�6��H�q"�� +��X9�����Q��R#�u��[�Pq�t�=��WPZ,������ជ� i����Mpn�C�,5���LL)�W)�g��2Fa�O��`��s�����^�JϽ|�%VgG�v���e��l*�*���gUH��)ݺv[���NZ�x���H���C�똆3y��J�R5�`.�=8����"��������^�Xs-�R�&���� �>s��h%U���ʠ��|�I��[ΊZ��iդ{�S�(� p�5�p��v�軺�I�-�ձb�u C��`~�u�!�Hf��Ր7�|����`��`)h)������g6�M�#j+�]�6���7�W*�
QڞD���%OkdiU�C�v�,rD����ōz��^��U( ��Ts�(��;~��|��_��a���)Ѫ����0�bI� 3T��F�����<�%��0���N�Uy�	;�H�4��R��U���.1lly噻�C�%�x����m���g��W�{�C�uW��p�O��
t���4��ƠG��V�PT3djEy�>��Q0��4^�x�H�%�#׫��i}R�0~s.I��qk�ڒڬ����8
~n�	��\`����h+)��ڭ���au�Lof�.�k��o�(Z���ɦ/(i����W�Hْg�LA�Є�{I7�2h�+o���j��!�]��3�m����-ˁCSVd|�(-H�5$�,�ݮ%埁"���X�	9P8ޅ�:KO����Bp���O�W�A4�hZ#PU���yV�V���C~�#o�+�2%ʿ�gn�_6�x�9��#\�#k�&�	�T���h�l���s��:�Y�h���Ol\g̓^!�{�<ğR�՟p��0ZY�X[��g����*�q�p�j�l��R�n%t[.����-v��c�h��԰�I\*'Y�[4���-�k�K�z�e���V� �b�v<dN@��;5�6�}�*eU����ךt��+mz��6#�qd[<$��"K��u���I�]�:��a~U�4�	�����7�Gq�%�����[e���͈]V��D��'}���
H��.y��#��W�
�����0���b�Y�/��1��x��I�@|�9�U;s����T�%��Gm�^�iB��O�4�8�6h�>�5�w�pB��온�������SLK,�K"�ts Ws�hY8�r.�zt=�@EFI_QH켎�h�nx��GA>X�w�1 >7g8ɩJ�F�1(�a|T�����﯀��;!�PL�r�Y��]�|냹}%��D��"�,K����ۂ���g�C����t)9��xѓw\%D�362�(�y�B��i&��4T�%;��L�����N�ʷ,e�.Ndl|��K
<w�=��p!W.(��e�xߪ=3����fRZ���{p�R0#0뙨!�ޣ ��!j��PP-���oEX��Rz�ݓq%>�[)#d]�*<J�*=�:Gr67jo4FR�	�f:������9jk�%(l0m�߂Z�Ǭ�A*�F_I���ET�7�?/q|����A-s
����p���	��J2��bih�E��NU�Zrؗ�d;����J����s	�v�w�js)1y5NO�me�6\�6���wL�Rj��z���K���ya�I�M�(Iy���԰���:�_���T�-@���O�wx�'(���1ۅ	G��R #�QR��5�놋]0��6�b)�]W0 ��W=%d��T��v�CM=�0)�%bl�*���D�a��"�fT�ƭB}g$H8�ݫ9ؔ�;���F�f�Z�8��>��]$0��v����E�0;P���K9��� �sCr9e�Nn�D�����e��Ƙ��(.\[`KO0�W���"ܻuth��x8�uT)2�5BS��"����U�0u�B� �O�$�ǘ63�o�ۡ�N���4X�W@O�o�g	3�ڵle�V�s���7�M����S�}���t��eV��Q�����j�dM�O���w���7s�aH���n��x�	Fzv�j|�np�G�������&!_����$��#��x��nt�ɫ�̸�wgv =���VtCK����7Ben�I�o�U0vb_�Oਉ4�h�e�R���Y3;6$�}��뱸�+��w��Վ�*B��mr��<{U0�n�{���o�I7Ky�,Q[H�J��C,]01Ĕ�y��~f��˦��0*7�\=ӛE١:I�%ǌ���pOݰ��}�ҽ̿..�d�9P�B�H������,(0$U�!����b� �k��M�1Y+����n�z�(�!���:��e�/D/v���AmO-�+��J�H�������]?�n(�~q��h���2م��z�8y�)�q$G`�d$�Wwn�I��G�*Lv0>�Bq�4ש'簓m���D&��6
��<��E��ȗ�������ǪaM����~�阒�"����[_�K������ĳ�c,��c����+����q��}Wϩ�sxG�p?D��4���,Eҽ!��A	�	�m@]K�3��
uY�=8�Ь�]��*����J&���̭���D�)�z�CW%���8���<m���m��(����Ğ�M�]�r���t}���PwB���M���.���$��u+�Jy��2t��o.�25�W]ᚇN{K=�J�GۥE7Iz�����>/	!jw<�v�9��@3|�↕aBC�-Ϛ�m�u�!�=�L��41��u**/#N�1�*g�M�?t��Ԭw��.��n��(~��`B:� H�������'}��A������J{u/V��ފ�w����F
� k��/�%	�-hAm?c��(�
�qm�.{ڭ9���)�dTm��Bo�.���6��L���P��I���j�>�MC�鿊���V�F'�^�L����H$^ipZŬT�0q��_0=��.jj��uX���-f5��q���G�y���ʺ��y�ԯ6�Ec�\)�\�XVE�j�C��I� ^RZ��(ͻ���2�[��'���t�t�J��G����ړ�ԗ���oA���7�?=��6�ԕ-'-��
�����'�6�w��8��0�: �z���$}���^�y��Rf-���,�G,�oƢ"ހ�2�8����x&-imݙ�Е4��;�S��GV�d��x�pB�1���/A�\������9]c�>&�#W̭*�;�_�O+$�/8�;�V٬��w�Ȋ��'y�v}�)W-��5d� ���w}Ű��[�c[��O�V�D��
�#�n
�x^�@�m���Z��7=� �O	���}#&_���զ)dڑ-"4W�r��A���c���pZ�V�y�>��qɌb�Y~jK��:K��B��L���m4�奕_~�t_8���,���KnO�亲�5R��}N����s�����O?K�n��>2x.���u/p.:�;c�������L�69��DN��|�?y�!�IݻyvK
Y�c��^nubn�@T�x���ܜ��H���&]����q�1�Fy%ݒ�0 Y_[e�#}�U���S�a�4ۗ`��G����,�ΰ��~�G���[��vhS�(|
��щ��P<%�~��2���Tgx�p��k�"���jw'�D�>����Ģ�5ç��( ��*\{8nC`W��
�}�����Lf��c=�vV����߉}x�$�� ۗ�2��~���e�.NE�Mq�N;�nwڒ���5��,�� �Ұc`=�[.p�r����d��_�ص�b0`�±M�7��%�C�P�ֻ��5z��#�&�Io��{j���|��� g�U����pR3����?����!Z�lVvc�~��M�+�A�X�D�f�L�5�F��L�&(l�cRkh�b4��Yѩ(����n��b  {����x#Ն`A�h~[?f|l3z�r��@�4bWn�Ha��QQ	�*�k��N���E���e���ueJ%э9��JK��@
�ߗvX"?��t������.����y��ɦ�!H�S�ƙ��1˰�������~"{�O�s],�]���NW��Ҳ'{�zxhr2[�	�G3�����5�v�f��{���ۗ��l+0(X8�p��^��	����>=��8�>�t"����D�n����e���.;�q���0Η�&�y���[���GE_,uߵ|��t����} ��na�����%�??gi$T6���4��̀<���a�䲂�p�q��m.������v9�qu7j��I��Sw}K_|_Y~���N��l8H�2�j[�F.�=�����@	�3Oup���V�b����>��u��@�fX��d���N"�� w�C���C�M��+��<�Q��zbb`=T�`��¥VE`)��&cH�<��Apb�1��t�V�0�̹�(B�|sX �3�s7����K̎Ъ��$U�,ސ�
R,�d�*g�y<�0ٮu"��� �0� *L�&؜HzS���볘#�	,r���6����3�WL�v=����Ĥ�y�5�F����	CP����X�ؠ����>7�����T����(�\*UnI�� x�����$$�|Y�s'P޽�����<� ���]��S�l\`�Fb��tK�G� VCb">ڮ-!�����^(�{�5<:��-Q���!jZ?���߂$�i�)<�O�h�Z�9���3����������2�ÿ�F�ew��v�q�*r����G]}2;���U(�B��3��U�l{R�hp�i�D�{�Vx�~���>����PpL�K|5���,� *"zI��X�����7�]١�l�D� D�b��7��Dۿ����3f�h�.�ٿ�'[��յ*_S�Fx�H5a�r~]#�&��1�<����:���S�j�r�@@�zǷ^�J�O/�@aĚ�|�~��*�Z~�j�4�
�*EvV�"%��ʩ�2�bu�C=�r$��l��JYB����7�[�o�p����FgD�:Ѻ���]!F�=�"�}�
�%P˩p�AxbA�h����6����w��8±�s���`q��l�)�5U�2T;B��l$�Õ����m2��`C$�����E��W^�88}tg�lX��L�t� �I���9�7�=ta@�Z�=��,��^g=@���|L(V�[��oV�-)��T�R;���@tX5��>x\[E �
�ֈ����C�MJ������񒾐Ӫ)P�9명4r�{�����&��B��q�bF*�(+��Lm�u�p	]�����r2zy{<}���דo�u
B=�L�՜҅�xՌ���⾌<%��s<�z [�Fɠn�d����<cR�(.k�|	����X����Y�(	Ól��o.�Uw���*��$�ҕGҿN���)���7��W����#�����6S	(1-�舋�Lbc���;�����e�}��-o�aB���&p�d��z�}vS���$l9�iܳ��)�{�e[LVۢD��`�hF����NrͿ�v��>d.J����U�~�zۙv1�ؠL��.�[n8{�B�%]Ԏ��wH�ʎ�?Ϋ���8���16��H.8�h�c�d��5�L��]��2���U�p�o��(���}!���iB�7X�t�jV-7���o�5��8�8-S柣��Y����3
�< ���l�^��C	E��M�'�Sd���j��Jxx�M;���C/m�{�*ɔ.�%!�0MT���ںi��4�
s�"G�̫��1�uB�rz�"dJy��R5�N���
���d=���S���$C'3n��x�x��z��}���t����G��F��F�^���\C�x?�����S�O))o�D4
�)s$D�����>OK*��|��O�սZ^�u�qmT_�}q��9(F�l��2��^e�o��xL9%����c|Ί�$�4R����>���	�j��n%)��/���ij��ƥ��f3��Z��c;+�攐8��ᑓ�ן-v��]�w���a#\�k�L�]�V�Q���u�8��H�t�0&������]7�.��UEݫ����v�FȀK"�r�o�����5 �_�و8�����n/�����)>
!^
�K� �6�D�Z6����TvP3ۡ�j�3�hF��3�L>;�N�Î�h��L����w��4N�6����ozq�U���XY�++�Ću���q����R��/*�M�#:�H�H�ː��Ʌ��y�ꄯ$F�R���X�Y��&�* J�D��m����wG���޺��Ws�xr���~	��weX�At���һ��_҃��n���������9l�ıO�e���Ǌ�e�em&Qe��bX?��ʹ�(�<�v��gRJ�dg{��y��ĺH��_�������i�?�a����m��Zh���	�����Iz M���г����� �K�7�v*^)Pb�����qu��*R�7��Je|�~����ܳ�vY�6�W:c� 8��,���$P��_x��3I.$O-��s]�F�����g\�Ⱥ�sr(�me��������٦cd�c?��n��S�G������AxŖ,k��(X��ںz��<�X�h��2	>���	I�Ƣ\��<R���XAy���T&G���e��A�����*B��D�͈I-����7p�6�O�r��5hO���cI�`-yW����T���F���;�.�[y��,�tm�!�)��8<���~�1�R�c�e�g;���H���.F�=���b��"��OI&�o\����40U�8oY�T�;���9�;e�/�⋿�2fϘ�E�$ҵ��d}�/�Du�ڞj5��?�Ѧj"�8�9��fo�^����Z2x#�L��}m��5�8>@S�p�:y��`���H����`�W�U�~�w*��/����y�T���K�o9" �Hv��^�=�u�X�fd��˷H��H9A��8��&��r��n <"��l2li:�G����}�	O�����p��a`��{k�
�tu�0f�޼��QA�ʝ������g�݆տ/��#�8bw¦���Rc��֮�8�W)&P�����8�M��B�����=���5�%�Ij�\����(KS��x\�˗�)�L��r�a��Q���k�؆BlG��+-���/����(q�����矆�"�l��� �O�eD��Ydt�R�U�1��R�/a����(�L}�2�=�;O�#"R�9iB��/����gD�tQ��
ؓ����O����q�Pr6��r�Ӓ�H�tj��%��?�r�Y7)��$��Ȍ�@��Ld� Z��݊�Ԅ}ʊ+,;N�	���#;����J�X�_'v,����N���ݖO�_u�ߏ�a:>�ƩA��a3���mJ5�;$u���K�H8+�-�z�}��?��jq�@�kl�U�����	R�P�.[�M��ڀ,.7�/#bݛ��w475��Y?�l��^Eh�����iƳo�=N�N��8TG�a����k����oӿ�A1�����4(G�`n��4�f'CZV��Y5��s��!ܯ�($�U��0��/1�|���-h��1�V��RܹTŽO���XO��b�$�lۘ�:���Z<ϢW*���/��Pr�0�T��O�Z���y��X�Z�(C]i�+�7��\d����iB��8�q�����������.�=r3����M�e0��T��p�;��tC���^�_����V�֋��p��A�hV�s��p5��`J�_01O~eG*�@a^ީm�`���ȈA\[Z�M=Iᖳ��4ߡ�?�ٳ��Fͯo���R��OS�b2p��"�CWi�M�4�(hc J�?�+p%�N��_L�"��N���|��-Kj�I��*T�D6�2��*C��j�N��wyS��iP)�dqPf�X���,o������
�	=c��$��.���w�H�׻�#��KXҬ��?�}�^�K@ԅ��(��q�wo�q��
 Մ�jN&�hn|��;���9�Fbzpsi��e�1��p��SHs��Î�͞�ɖ(��[�};O���,sL��y<��0@���<�v`��}L�a�f�o���C2���ׁ��YWn����[�iEM��%��mr��l7�7g��Ƭ�wm���CJڈS,�ַa�!����M2�5h���*��sy��v�E�	�ͼ�,)�5� ����S��s?5bǚ�w�+�[�tJ�1Y��{��3�Of�L�#R�x3Z�s�q_��f5F�\+L����E=�p�������.�_�����K���4�A!S���a�SkT�fV���%��V�H')�Ma8)��#0,1�Ƕt��i����ِpE�ڞE�]�I�R���ajx�ٓ�Wt�D�*Qjvz�H��[UvPm}�b�+�<R�����{��-!iL�u�2r\[� $�ƙIf������1���Ex{�<�+:l�ł����V�s��\*6��K�\��>y�vA�@cN��ǻļl������Ӝ���~�f��˵�kD�>f8�)P��K��g Vo^\k�������[�Q^�rt%�'�R��L�_h �Ē�q��]���j�3�Ge�/j{2G�l�dO0B">��铲��KҾ���:)=�Z�a4��;f�:�[����"����+�(sw:Q��BW]E��Y�٫-�z�t(l�m
BhG�e��Q�x)P�N�R��1���5�)Pcz Jdr�J@	��4i��4�J�kV�x���iu���>k��y�S�&,��v�+�y��\������*�Y��v�K��shɑ
b	y�E���Ɯ��W���#:%��)�4FQ�k|���nG|�]Vu�Դ��>g��/�]8������%�Dg�L]��}��l��r x�L�I�W�Œ�@��_��_�M�b��=v�-<����x�WGM৩��<��UE[\K�D��p��9(P�-�c;��#��3���d��XP�ܺ�vJe�\�3�S,�g�������|�I� Ks.m!�����(s��6Ł#����s�e��m'IrSל���3��Ŕ���}�2��9�xw-k���;_���^p� �Lh�spc���=�!���YAH�!c��EO�:"���)hr'�{=D]�)k@�$j�qi�ꏠ8�w�f<�Y�������	�8�C��d18����D�B��,���&x�o���ۘ�۬�1�7�>�9��4���T˴]��eU-�B;(P�dv����]&`�u���S�QV)T`�?�<�woC��)����p�}�)U3L��̔�Hy��8�� �ܕc�*� ���B�eȂ��x��Աh�<z��,w� ۭR�q��V��#U�*��j[�(�ԝ��.b�d.3�c�Qu�xT���;�r���kUr�o�I͖��C�3ܬ���	<�9���
�&�e}^s�I(~j��eP�����cy��1�+�M�����wg^u��"�\�|-��=�Q����R	l�d�x�OC�hA[¼<�!��HA)�A���#��8f�<B#���ӧe�b{"8T�2)qX]L�<1��3�'�r��R��²S�h=c����DL
��A}v���Q)e�a:'D�7q��C�ā���0]""�R�h,/ȡ�&G;x(�~�|<����W�?��ɪ{3,68ci��Aik���0�m�͵9>��P"���o����A����3�㸖op:� �LFc�b	+-���-�"�ױ�2m�C���O7R!8�H�HV5�26t��RΎ ��Tu�` ����U͖��6x�I��4c��@YV;�7���rG�ʌay���/?�s�����T�;�������m�!���`��n;]o�O�C�2q�ɴ(ѓ W"�ЂYh5dl�u�f�ϓ���frv�&Ck��&n���B�U:�Up(��~Pt=u���16X5��=s@�ym�W��R+�m�8��'�伾�5�q5��w���1;Cd@�#�5��;֜2�K���� 5���s3iQ���!�$a�8�\�^Ыi����=Zw-�_��8[+�j��Y����+햤 \��q	�v���'�t߸�_�p6���S��L)j�����j���I���[[g��Di�ͭa����jh���6��U��RY�tR�{j?l�M��Ե����~����RR3t���$��Ó '���Y<���4)��!@X��%�a������U�INY��:��z ��-"Z��x��,��(r �w��0�_��A�01�p����a�߂�@��  ��Jmݟ?gAU�2�D�O��fוҾ%KX�J�c�I�	.2��^I?��w�B�q��'�{[^�ҁ�qެ�/rHS����Ր�GZk���}v�����\Dc>9��8�;t#r����C!K=cN(�XY)_����iL�[�������,O�2þH5h�i�SYw;[W�f��V-ͮt/3Ųk�{�(��I)F�i���^�h7��b`q%��L�Hg�PDVh
��~�J�<TQ+ʗ$Y/�$�����hl]��@���?e�z*�k�]ջ���dNE	C��.�#������S<`T��Eķ{�5n��{�N�T�4y���S�����u��[/�xc�rCKH��8p�-��c�M�A,=�ιe��Vk�~F~E�}��ь
a�m�ʒ���T�zh� )B�,Z�W��5�FF��,*�b(�8������2H�"X����%�h�u��6�ft�q�O��o���b�[��N����T�W-�(�n<�Y�ez0t��f����j��[�k�r��	�CDJ�,�$U�_�q��)g,=�\���Ն�7m��5?h�l��k�0�x����M���&�T�Մm��+�蕵@!w�HNx�}���0膯ew�Չ����(��X��G�g6ZDZ�D2�gGWϛ[����a�e0����jBJE����%8D���Q����L?�j4=�95${��jg��yaV�V`|�$-1k@ƈ�A'
M�D��u��w&�JՍ�H��)j��|�Ds�,)��i^���B2B��ݙ�˚E�^�\zyT�-ҹ?��Y^�(_�'ɦr�+�+N{���8�<i��ud+]5����'3~_���6E{�՘�����5�w$��GP��0���C���[?���~��*�{ֹpO�����cU����:�E��ع�qh1�Z��gܰ�	�}}[���pJ�^��b%>b?��:pL��Б�a:��>-�/OB(^�/,.c�غd3�z��p���[q�-��rN*���i�E�By�?�1�{BW�&��b�Lޡ��=�쿣��l�xY�鮆����u���Ȩ��Q*Y^�V���B��y������C�0hJ��tβt<����l[���?�8�I�ʩB��Xl�8�8���V���a_ĳ�j��{� �-����Yu�vH� �P�	c���5����T�"��It���v���o��l�2c�q��T*�G�nqt�@�8Um�6 `��/�f����1mڧ����WƘ�/������D����Ƽ�>��1S#�cI^��~��Ϛ��)5�r��ƹba���?�V2(�1�6I��A�aQ����ڰ�:�n�=w�����KPh�i״��3S���5v?�w Udo����������=`�8��s�У��+������_�QA�yG��.S�L��>�˖H�G�[Q�7�RoGu�n���n=[7�$��s�r���.Y�������K��	G���;_���թ�+q����@~L)TMb�����4�ީ���7B�e8�c�n��hL�u �d�]R���MoT���^������\�r騧i�b&���m�z�EF�F}�_�.C|3�c��&LT��v8�����9�;ވ���o6vKЀg|&�s����7:̯���*f0��:���l�a8��cr�ĀSB2����:�<�>.���d�n"�&��{>n�P'������7��;P`��9B7Lg'����L_Ҳ���$��`�zr�v���M�(�&�G�)����U���Z�٪7�z��|=�ͽ+�96 :�����!m����Xq���޺�]R%&��j�4�֣�� X�p������ɔ��� ȻF�j�u�47h��Q�ֈ���-�����ߟWb+��״v�έ̠j�SPVgP����;�I̻��G?�=���z)Y(پz�����GܱuR �_�g?���1��W�g�����Ǯ�|<�)�o�x��F�z-�ٜ�4g�Vf܊�4ǍOQ8C;4�a�/��Yt9�֏����E����l�
Lb.5d��U�PR��
�J���;����͕�Z80�?��=���ߐ�3�qH2���?F�5�]��H&�S�n@�YT!SyFk��'ɥ�L����b3o���q��+p��z�T�^\Қ�O:���Hx�-컶e��H��u�|������`��'wH��i��o�9N	��ꡝ�����v�*���;�;6-Fm�[e�n�]^�(Á�WEG�� ��������~�|zv�<ϯuyd��6P5�H�$�:�����R/:gB�,�j��������(�*tj(��KjI�c
(S��e*��C5�7pD,���{�u{�
}�����Ґ�$P�)�<D��òF �)��|mN�����k�>�	���|�4*ڭ������a�(���ݽ��sD�?٤�lN4N�W@��K�OCV/f>l57�G��^�+k�+p����t�AOhp�`�S������3J��G�ɯ�O�%����f�@�x��	x+��X��|�4��@�+�����s�˪G�)�ͺ!���:�u�6�]��r��:���+#	��N(�11�hA?�eWPX�l����H�;�1z�[�x=�p�@ۘ�G�~O'�?�C#�� s�-���6=��5E�dxJ*:�u��([��� �2����Om@׮C�d��gGJ�O�S����I:C$��TF���E:�K�ó�����9��5y�J��5WI;;jϺ�ٹ��Q"�uTǬ����Fq��[�F����W(�+}P�Mɾ]e��� %-��:���%����/Ki
��m�G�e@�>�������T��!�n�O-�yh���̸�1�u��rBq�Bf��@)2��7� :[��O�Os��T����@ �J�U3�z�0��.�x{�|��A�;�3�}s=�v�9�XRc�tc�e)B�I�vȶ�WL��70u�B�����I�p��g�����+9"Y��+-�r�eIp
��)��z�HN�`�oѧ0TW��c>�sX���o�,�"|AYrJ���|�C'��`c��eت�ֈ?�yj���ya�4�����q�x�-<�pÔP����d;#�pҘ�h;&ә0�@����4��eݹ��md^��2�a�]�����KI�<����Š�	s��Rj���G��R�sz���1���1�4
�%,��1�e��#o�X�H��d���|��T)���]���c#���_[�	}#ƭh�,B�{����^ �yL�����X�Ֆ]o�'gZn�٘a+6���3j�M���Ӥ� 
pP����r ��{���{�"'÷X{c�J%�9�����*�j�7'�/��c����1P ��\�0�V/���4��Uj0ˇ�nJ�T�m��y�`i:#&��=�y� oyU�<���j���\@�{(��ܒ$nE���]��'�����q�<���`�G	��L�Q��|`��!TBV�L�J����`LA�kWd3���A��'$��O���d�,��1���%w�B�Ϭ'�����g���;��
�R
$K�%�+�G</r�~A	�We�g 7a�d{f{t�B���Sg�̖<���1����5[yv80j\S�9HuOs�U�;�l]���:pХC���ŷJ�]�E�V0�̗�@��|b3��*�s����n�L�����V{X{��%�ۓ���K`�SR�m�*�ՐXP�M#��{�9`�笓K���cK�9n�B�1�� �(\�ؤ�� Z=�az�+H��erd���ըI�751Z��mN�ʁ�~	�K�z��^���RCi����,E�}��j0��?v �ځ2��mIJ�
2f��o������׬�"���jHaG�>����8%g��k���r2�ᛁUݱ%�'ۘ��"�E3g%�����j^���q�S��BvD�Щ�8S�����]`�c�OHi{�}w��� w�-k��iJB��%U�9�{�X���d'��l�[�RR�����9���ܚl��H�[�􀖎�!t^��ztF������ж��
q�׆!�ԫ:M:���D|��]��1r��p3ȫ�ףJ��v��y����@���ۦ5�$����ܯ:ji�^�~Qp��=s,�E��
Ϝ;��G�][��ȅ�A��Q�w%YQ��f��,�)}==���ˣ�D��ټe@C�R?�@����9�����IX�V���3*��Kx�@7�bm����( $ �9p�,!A�k��8�jQ�V�W��!p��J���U�C$W���2�my�O(C��,:h�3��G���tϭ���'Ⅲ~�C��B�6���ޫ�r��|`��U�qM��^�nG`��)W�r���^���?/k��q�7A\I���	�O��0�R�y��N����i��-��g�(ȑ��m��n�t�;L@�Ԏ���H��2��t�e�B��U���&E�oev1���f�lg�R���m�iă6��Z�,߅ċq�Y�����iĵ�m �����$	d�(�4��.�"��>���?�Ŵ��Zߺ�F-wMKkטȕ�ȳZ��:����PϠ�R�?��N��%��0�0���ԆQ�~�wx��<�ఙ^���@ʃ҃�dj{6dHiˊo]��f�3����h�JL�'��^
:���H��]���%�j2�ɂh-��xE�ŧ9V�n#�.�3g��% F���&��h�#����v�:�ER!�C:��4rP%'�KH癑|��e�͎��(��S�>(�Z9���(���_����t��Bx���uH!��.lW�d�,.�����s)˶�R+p��N֌�{~{�!t�O��z5. �9YW�a�AogYO8jF�5G3�CR3"�T�l�Fr帜YF̍neA�CE�b��aY�MJV�)wN�{�r'?:��6�|[��H�|��'O\P�Ct�5Zm�R��ٻ�Ə�8uA�ͦ��/k9J���Э ߪ����!1��/{
 �XIRnĕ�3mcՅ�jw�����ݩ��+��c-�8Am\�����?\:ӏN�\l}1��t�k��bi��
ܸ�"�!a(�b' �ը�s���_w>u��P~�k�N�;f�q�e �CHC�&�f@O+�@���A�U��Z���{�P���N"J��J5oY�����сvC9c����<	�\�8�-���Nv��&�֐%g�1՜DR�N̹O�3�����:�:�K�	ޔR���?�,��j�X������"����d� �j&�cT{�܍��H�m����Rl3���戩�oF���� 5���w]C���:'P3,���)[���J*cz�-����bbi�V������@+6��Zp��b�Cd���߷�4]��l�?�vN��yW���GpKhBf]C'.�VlYJ��r_gi>"BV�F-Ӹ��}���祼�\�?Z��h[u�4�L|��{Nր�&���n��U�Ə?��D|�	<���Q:��Z�4^潔ı���c�I��Ci�h?j;���hL)4�D]���Z>8y��!kT9G	����x6���*�a�k}
Pca��k��,���&�I.�)���m�D������s�=���-G�?u�1�*Ƣ�����H��w�O���yj4�"�^��Л������ז4���ZKΫ�A9F��Dc5m��rǧ����<8�HD�B��~i�\A�+�Z#`���gӱ-LE:�a}�Em0��p��ENP3BCR9Hի�z���h�L�+ȫ�G_�Tf�b'r�a��bL��$�vc@ӫ�L��̖�	v�1m���\���C���w�3�0���G:ϖ�ާ����4t{���%����!�u���D~M����Ja	_��TqN����j8F�i1m|ܣ�O�y�YƖ�����ptjo��n��ٻ��7���o}ǡ�XXӅR�uMa`nߦ�H�=��0�ۭ�Y���b+f�$�g���N�g�]vl�����fܖc�E,;�������ݼ��_c�l>kw�;^H�utQ���N��`�
�_= �#`+Q�5l�]����t�����'��n��9"d�v@����X��j��@8�<S��Yd.���z�<C��O�Q�6�4�� �z�Կ����p��Rq�Fkv��VE,k��sC�g��6���(�h�U�+�T6o�ȡ>�̍Ķ�Le3fՃ���-m��i���p�s�.�%��X�e-��[��P�[��Y��kz�y}�n��n'�4K�F1�ό_��~/�4.�$Յ���1����������lφ�5ƹ�V#�@�Z�؎fUS����%a|��E�@��΢[���yg���b���ԁT %,�C+α�m 1���Ɩ	FB��hVR������ ���F��r�7;hƪ�ߤt�fRU�ܣ[G�Iy���~3��<_�#q)��~xh��������Œg6�q�럁�Ӄ��#���;���p�4����ܜF9;��
?'�K׫Q�4��ȡh#���J����
z~c�(��y�t3I�$x@�I@u0��"��^�	��QI�?}�d?��I_���+��"~Þ��i�� }P��am2@�e��j"��YJJr�,\*��Z��_K޾�C�Z��?�jn`=A�C�a	W�T�/�{����h:���w#��ZВe��c�#� �!��쌈��	���n����j'��=�0��(6\m���Ho���\��x�il>*�[��}��Q�+1�L!L�8�s��e܉�gz���,ӡ�7dn�FO��kIG_��>{���ҙ���h�r�G|�C�!�C"��=��B��5� ��`(�K�?>X)R*H����o�w���ź���.���Q��d�ձMJC	@l��q]q���|��8�7D��`%B���FL�t���?��%��`�TD�1�d����>��I`�����΍�(�v���k� pӶ27�Sh�b[����1^�_a���r�PG�����?�6��9@U79Wf@��{O��F�بa�0w�{	�k2�̱Sa-p����W�
mAU��3�G��(p?���Z,j��z�,���%1۳�cS��9���;8��R��\Ds�Dn���M4ˁ�����e����ˇO_7��	mD"��4�x���xW�C<���XQ��|�W[#����Ğ}t�y�V�tٟ
���pM�4CKi�a�d�t��*��J/5Ӈ�lǾ$�����d���]`�����u?e��E�|�_�I��F���eӟ����y���I�o6������)K�OB�<:���*�w�L�'�xN&�Ƴ.��WF������� I.���[�����
5Z��|uJ��w�H�bYш�A�$^oK@�F��ཤ��Ǔ���
N��b��<�\l.��}����F%K0����i�1̸�@���I�-�S���	{��9��O�0:ɑ�Mi�cnA#��h0���x=V��vF�vD�rV?�>�ʚa�֍ �pF������N g�g�c�Y�'��h�MwN+�����-�naJg�a����,+�|�MPB��;�ض���Q�k*ť�+�N�Ae�{P��3n��oZc7��6J 5t�� ���w��_߅u}{�U�?0�N���M��Nye�I0`w^i�����a��n�Bv�m���Q-)]/4NH+3,����m``��p��";�-�P��B�;�%�J�*���J?�m���20ZR�c}��۲��P��q���/#kR�N(�͏�[1`������m�OSŢ'F�R�
��ut���@�5ܟ���F��3e�.�wD)�q�jU��C!7��"<ߵ=���s$���T��5������2���yƷ��e*�R-�-#E�%��Fc�U(�s �7�_�z��8��IA����9�QP��A���"���u�`:ugI�4�Όc�oڤ������D}���P6B].�ӛQ@�R������þF3[!!�V��.+�DUH=HӦ<G��A�\�?�	�G��E˻M�xɨ���I(i�C��^ IP�i�fd������%od@��r˕���Q��Fa��,�J�B��1KX7ה����ݴ��=Wz +��WA+7��������!��V#@Ys�s�R[�]@�fM!#̦�5�
����6�*4͘}�k$�����7���_E���	z=��Gq8J�t��C~�9�������Y?&e�LC�Cۜ�XQ��Z���.��Z�t� n�:�'���
ˏ���]Q����V�������%�ka��HQ������5sRz���9�J3e�2��f3�楲ouz�ظ�t���^��P)9cb-+��:h�c�q[ONY.+�1�x۳�5Cъz�"o-�&r�*�x�xI�{6^xM;!(4^<1�����f���rX�z�� SζXZD����}x��jnB�o�c�k��t��X�� �4E����o��Ig�u��]`���6�CbO���+��x�k_̊w�F��e�a*��������Bݝє�~*e�0�'�ť@�'����8�ɚ`n�(-��y�]�V�i��R��svs�9k ��K�+����+9==�������>����r֙Rma��H퉦�B�hj^��>�y�86D9�pCbD��^ ����0,��:�rAl�5��lD�el�������\�P3M����=p�/��x���v��X_��E��J�ە���i�˹��#>�N�'���ْ2Ç�1�"�_	�[�c��"[z�d���1���W�Z����jR��f�F�Bo��Jؗf,^yd�.�����۞��aB̌��Z�_��s� �K��� ���)�V�B��+#�y���2=��	)���ݨ첍"� ��nƃ���z�Ao��%H��ºw �(��K1$�5{뙃�ޤ
E�����)v�5����N�pr��M۵�N��+�@����s�!�C3Y h��f�Jy��Oʖ���쇖Y�tA�iL���I���r}���[���9����E��=�Ώ��aݧ�����k8j+�l#�o,�,�cș���c���2�F�g�������!�h�� �}�/�1M��{�V�ٍ}W����*�%�H*�QJ�,���gv|�=C�7������^��Z�t�-��*oK�E�9�@2���U�2���5C�8���%��Κ�p ��QV�	�Upe�3ZBA��d���WܻdFh9Bh�WiU�ռRѮ6̏��aԐ<sK����Y0�lMz���(�jK$����)u�^?9�8�<I�}y������Q�ۃcBKo��7�P]�B�J���^��}�$p�FDG�<f��{�����iP�Ӏ7�D#i�[�&�F�ȓ�l�٧c�d-��&s�;`�g����PV�@|�
\蝾Pl��c9�(Y3K������V�2��؍w����C�I+�m,����g�,%�l�@ �k��~Qo�3�X�'�PG�f&��RYj��w�W[��D�-�����>���q~�Z�!�'�nPd��5�����\㧗I��l�=��TF�����(�[a�����w�N�1���Ӹdl�Z./�񛦉�=�^[�p"Y��wޗZpy_s"�@�T�ցO��B�#z�A��1ʔ͜��u�q��|Q"��*@>���Q�:;����^U`�E76�St�m��pӲ�zѿ&2x�[:�-��!�G��^W���,���&2C��XЙ�4��,�ؾ˪�O�F����0!v�����!v4��������$�a��1H-e{o�	��L���m� JGu��s��/|�-��m��J�%�L?\`�Y�b�gv���+(��l~�����sTn�(���i�R�Cám-�(ɲ`J	�˥�_(9��%x|� rA#�1�eiv���(��홡�I%����������d.��!C��Q��;,y���u�9"^�СX�]��<l�0eN|�̬?m�Qy7^�_����o�@�U�o�Z�q�c���*�<4��;"saԶ5�tr�FY�P4y�ز=bl�F����z�:�`�F�*�؀����������ƥXLq��UT��W<�5s�rt� ��uvvG�z��~�؆�h<��$��*[(pǛY���/0j�S@����w$tƷ�ΥP�$Śe�	����*��6p��F��@�� R女�
MqG�	Ow�w�h�B WFO�~u#�Y�D{��\�ź���j�sf,Q�����U?�2�}4�4e�]�׷�6����T2����b�����w�o����X �IE�9��a�51D�Å�)M�4(�j�t�c�*@n���#f�Y�2i?��͓��i7�����
�~��"�]���z����u[ςV{�H���Z3��E�o}�r��Հ
�siXk�	"r�c{)����Z��j<��d����:�e)H9S���*������M�&�<K���q#wⰭ��`m�Λ��NI`���h��[�%Kϝ��/�
|��K��i\����Hu�y�Ŭ=h*K2f� W��������sh.����$c�!�p4+'�4}x���w[�|Z@]˙!�w����şCH���0�'�A���y'��^\��C�� "��;g��r���k��������R�Z���
%���S��Os~��2I�`���̥d���ᏏQ�hD~XO��F x��:�_F2��:�~7ӴD,0��жMŝ"㮌2�-�$�̄R8�\��gc�é�a%��!=<�5v����oV�e�	�{�b!6-9q!�!u�/(	_S����Z���қ���k��3���á6c�v��W3�b�ѽ(��<4�:��$n����\�fY�S)���+/�GLE\q��̦���)5��8k���y�r
� É��Xؤ9.	��E��"����Wt�j�2��w8J�0��33��%�G8��D"�Ο#,ϯ�i�����1��+� ��B Ʉ����{%���R�_M�Cl8�a��e��,��s��yK�ٛާt=�y��DP���N9angS��	�^�e�"ס��6u��F.Z�1fȸ��hq)[�g��-g���K20�U��S�nr{%�i�D�L�>U�� ���1�Ơ�/��I�Izv�����#cؚ�sƥu�q�Gz����?��/��f�!�sPЎm��ْ�&/��f����KO}��܌�kz�p�S�О�ۇ1s�26��R��L�=.�,��:qP�b��K�J���+^L�6�g���Mr�&�������<�FU��X��+�C<�S*�8\���%��"@���R���uC������NM�-l��l9�e��ͼ�_36�	j�WX���jkgx�����9&�H7�=�0� ~4KX5�����;�Sn�U�9oS���Np�=!�����a.�"�A:$�˨�D�B�`��e��Ygp�?���K�"�;�جj��m�R��r&rRQP��q1IZ��Z����2*=��Z Q�Ն+�K����x��i���π��&�r�C*j�+�b�p�\��߻{��$�H�D1$Q��s�a�J�*�TA��VA�d�w�sZZ� �����ŀRJ�쏞@����_h�]S3��5�� ��l�������8gu��c~���z�����B��U�����C��sI�����q�����j�?B�l����!'����5>�:h�啧��%[9k+|�雷`�%��]���)P�R�����'�h2��q�[�̮�"U�p��t�?�@�#�-"h1	���н�x	2/6��v�ړ�Ew�6Xή4�*6�G82�5̛V�vkt&)'` `6Iln����S�����ͩ9~q<Y��EH-�M�DRR����P���'���3Ο�q>��@���w�5:������;�	�	��GW���J�I}��].�(ý	�K(_�޹�kT�"È�#�r5��>���I�ȯk�th�Wʤ&멷	�D�> 2qى��x�m�IbG����7������a"��竽S�2[��?�X��Nk[O�3�BM�m�� Ş�|���M��0݃��laz����m	6���K@�'�Z� :�En��0򧂝�65��@��� 6A��Wg���*4li���_3��my���%_�h�#�y��|�w�LR�r�7��%f������H��p�}�L�n���X�nӔC!FO���s�<&4�8��E���SFxa#�<�p;�ښ;Z�^��ŗ�ΐ��	�H�����cc������O�Hr���F����XL��M|�Dh�qn����&}J":����|i�#�R�QkfD��p]ޟ[DR�mT��)���\�9��̈́X���l�Mq��$ ��3�����"z��x�a��嫌MϫNu\�u�V�]��BG���[[K��L��5]�)���\�����ewQa���1b���N�3�B�r%�*�hQ��z�B�]�&8��O�C��['�7�E�'wt֋�L��Vab�4�0R�3�$m��}e���d���%^c��[y;�@U	)��C����)����O�Q�<���v3��(�A��AjJ���1�	�|g(j-�1�n��Љ�%�����������s�8��N<��p��׌M��VEa�#ESR�6����m�]NF��a-O���fm�J���
�z�m��'Bkb�io0�/'�����&L�f��I%aA�J����q��o3��\P�m��	�v���l!`��.�c�U!�/��E����Y�4�Y��~��\崽A���&5T�[��G	w�p��J�w�bZ�y�=�aUCɽ�r�\������ �良x@���z(E���/�8�)Fy*a{z��ߌt�!�&�O���;���|�&��	�ע�:����0�t�M+�Q��%u����j���_�3+d��ڒb'���<i�	�L��u�7�P�G�j�H+�+�*l��݇�݈�z��]NHE-�|�/$�`�4�+���-#�ֈp�/��7�	c��c%6��]�C���!��_���1�9 	AC2��3�i��TQɝEy�-<.塯�l��F-|p���ivq	&��<s��z7������������i�NeRv&�>S�q��Z�Ot?z��Atf��T��t-&��8�c����N�|R����?��1����4*�m9����8Ʈ�"�O�2&��_�c��覑�>@��Q��kr#��18�O�1H�� ��;"��F��Zfʹ"p��$bj�*s���L�H�{�g��Qť�����V!�7�A��5���!��N��s&6/�w3Õ�w����N5��Q�j�V��%�t����h�F�%���y�\���e0����|�����ހ*��Ђ"8�?N_�/;إ|FESz�@�+�b�K���q(.�]U����6�9����1o-#�Ahb�{�`<�u)aw�RFj/�#�����!�n��}�jh �gg����V����XS�z�\�	8�TՓ����7�'���r�l�}�du��p��y�7�`�*M0Ƒ����?�9h����!2&��C]�������������h4��Yh�*���}q�5�Xhu�)�o��Ac 4P���\kpv�P�|i������ +D�;҂�;�9K �j�g�]�LW�%t��L��ð����4��#$�9�,� 71,��ݞ��n��|Ͳ���Ek,<��a� nST![�=8ϛ�v�%{5��Y\�H�D��"���$;&�m�����ua����e�w������������PbI�RlS�&��$�	RKd�ﭵ���)�o��>:^��݆đ�6L�?3T@ǜ���X��J�_>NV-�?��_�\M�����Bs
���5��4��A83օ7A���FLpf7E�����g�÷�35h��yl�����6^�����zf�K�]�F���/�HR�ݶ��n_�sw�w��E�ڋ��YK>X�5����=��n5��Ӫ��2^p��R�؆s�p�o�e�	P�+Lyr�¦���l\���X��L�z��]D�.vb��`�yk2���tl�p��/Ts\a�Ӧ�� -���LO�!���|���ߟ�<Y�~�����>��]�ʚF
��C>�C��5Z�4(Ȫ����N	�	�Smn�A���s��V[`����6+��C1{obiZ�N�)!S�砙�����:�M��v7��*K�j\��V�/�R�ǽMi<g�S���4|�t��[/�G�2�q���&���F_�|���g���r!�u^K�֝-~Q������4!N�_,I�V	Vkm�{���c=a|�\�'��>b�H��C�a��>�U����6�h��e�0]ײE�h��ƸD����p���}��Ę?�G�.[��"�K���2���mlڳ��Q�"� ��g�[��,�QΫ�;7�О_�!U�MK<���w��it�C�@0xa�\>��-��E}�g����ҏY|��V�Fn����m��vIn,��M�= y���f^�O�k�=������/�^���_�U��,�^	�9�C(�F����IT{�����S����i�����n�>��+N3f;���N��.�^���;����Z'�]�Jci��on4�3|۵�4C�1����}��GJ����d	��lk�0��������c�&}(��S@�=5�������ס��U ��P�Y�/��e
���1XZ)�G9�/����6�Rrw{�P�Y06Z��[�{g�Kr��΋B�|z�uM?�9�v���'��WŔ����ǌ�f�)�n���]�����%\�/-mo�,;��p�3vǺ����b8jr's��()![ИH�s���a:7�}�'�D 3d[%i������1W�+�z-��0(��^ZA�3���V��*�xB7w��vX�k��ji�2v����<#O)��~��co,i $���5"��}'>�rx�MpIpi�|9�s�O{��J�;I>FY��~ܤ��$��?#�:rd� S��	�5>����R�S�P@W(�6��k���әM�xm�+w��y��!t��*o��������SF������uYq�i�j��a#�Շ�\�1'���Ɇ�7�$�4^���K�,rW<��-�&��S�cg�l�Uk�^;�B����n^$����o�Kj��"� �K~�X��s�!i]f�ȤX��S���D3Q�����(PZ�����X��>�m�b2��p�C�.��e��B�;�,���������g{��K)���ĺ$cݰ���(.f�cQk�tǘ��:��e��Β�w�Q)60�v��O��������A�*�tڡ���j�F.�K�TU���06]s��ӭ��[�}��S2V��������^���`��emsm|PDq�ő����^@Έ���h���&I��cv��TT4b)_���U��o%c�K���m����?U�go��7����E�f��8���@z�\�� �5�����
n��vF�!@�ܪu�*@��9{� ��&�v-)�� �TK��O1�ވ&��+[Ot͂���r�)v��@��d���V��ǳ��t�Dj`�������z��i��U���d�~·�L?��Ɛ������MʢY�@T�s�!�������;��j�� %�E�!�����d~݈�I=H҈^H\+�ɋ��*e�Y��/�x�y�D/-�ϾOev����o���V����Rwn��`cy?\�\���w��]�0�5�������҃�:���Z.&�qG:���q<���48�SX�-Oo�T8| `�({�gs�����v�e�z�����A�M@?�AjϪD����3#Y���I����b�9"�ͳ�؄��aTM���#Y�ݪ>�v�R͌YS*%p'۲��i��i�lN��i�٨*�x��������L�J�����S���
ַ��)�OM�;��H������l��Cgo�6��#��Ȯ��N����:��� W|�=7�#L��_z®N\m�Q�uR�'�@jwg���%��~b��[Os��]m������񏨢�(�bo�WaՓV�J2IΗ��ҭ=�ߌ��� �ˠ_>y(XR��0j�1���2ֆz�W�Th҄�:4�g�g ��+;��0x����T��1�&�8�=�9��m��X������],�q��ͩ�
]F$��j�̴�a��Np�%6��TX�n*snt��>%ץ���PP�@O���Q�\l�k8����	Bk�Š�Y8�ď�x��cd���Y�6�R���bc�	(�[ZY=����:��SP�s$��|�8��{b�������Bk�]���ҹ|�r����!Jv�pM'807D	oCE�A���
]a�w$�0d�5Ŕ�X�~�M,tSI"ѱ1CR$a�ď!��u�)-���Z(����e���%[)au� ��Fi�!�d6`���r���W�3b�+�h�D�:A�^�Y�d𯇃�̞�V8�Ìv��M� cr�-�E����gcþ�m��5�.��]u���-����K�#�Ԛ�g,��T<Pz��j��â.4�&�Y28\��z�ig�k!������Gi��p��!S=§�n�v���~c�͖.V�=lA�F�0N�p�*,��z�"����cAw!s�v�,LV�ռd����8�V�/��s"F�>	a����'<8�
���>�q陶�=y����C�9N����E*d],#�@.�8��Q��vC&��D�Ə���h?A�F=뺏�}���"l-�gIT��tn�_J?D�(Y�\��P�C�U���.5|ϐ��e9@&v�I�wk�����B�d#��/Ą`���*��t⎸��q�B��) �>�%�:Y��#��{8�ap���SL�P�!�	~;j�R�İ �a����i��wS�6{�W!��t̩	Y'O�<%3�\S辳���V$?��,I+�lQR ��o����҅脤�eq�g�57�Uɵ��I���Q4q�S8Ւs��M�����|]�v�0�r�����>�BSX��gPˤ��fȻ��+ǵ������45��Z_W��r��A�|k� �E������-��x�����`����ŏ���~'�6WǴ�Q�m5pL��t6�
�5� �~O�sqM���4����T���x;v�,������a+�U�M�B/^-A��,Ϻ��� �Kg����8��M�˺]�4B'j��R-��o��vh��J�'��,:��-�޹�*��I}��CV������'s]2�xt�;a�����N�p2n�Ά{�����D��܁��P=�*�F��޵�UI���:�i����#h��wʹ�q�6����t/�����v��E����L,!�f+uYF�"G�F^��ZH�"X�[n�y���(�jMt�l��.!u�z��9%��}8$��%.�8���嗶HB��?�尊��f�����ޔ� �Lݒ�~(�,��Q��1��}Ma9v�R���NK����b"ow��(U�2�<���K�V��_��V�Z��&+��E��,+�k�ܬ��/O�ꋉ��z��\�����R��h�.�MFb}����A��<q�􉏽a��������Ä��S�R
�R��4�4\�����n�l@D�xFC�Rg�x���9�}s�����G��^����]����7��ߙ�;��(��b�����a��R)�������ب�z��8�'D"�ӷϾ�b�lF��+rM��ѿ��#C<��'�s�O���N�g\X-��h!XT}�T�S�@Ǉcl(��g�8�媸2���E˱A�9�)c���`��˻�G��5W�9��Qaݿ/���h�}�ifXlF�V��)�Rd؏�~�Y�S&���d>?E���%��[9�9*�Ұǡ>�4�k����z$�*��r7{�D魻���[Z�u+�O���Iu*c`��#�1T�6F����_z�,�_�o��7	RF��F+/ia҆���ǟF���8|u�vO�k�;����ʟ���}U����O|A>���$�f�v�R���Z��������ωq�8��A���~��.�<��(}�Zi���giG�0;sY��y�B9HS� w0,�u���Oa�Z��b*�GA#~,@�pv�eО���f��=.8�C�ڡk�̀�1Y|�ܘ�������u����������c�I�� ��H����m�ÆhFf�@��.C�ڝ�|"�E6v0��y�Q�n�E'�L�a=��t��Y�%M�i�^�z$�"������BE��*��~�n�^ ���W�����F���˟H�><�bs��=��y'�ȧ�_���0�<�X5�f�1�p	sa!>ѕ�s�i�	I���ۊU��Cm @0י�.�d��ü�fI�鲊��|����e��\������	qC:`1~vò��J@f��Wr��:��k�o���Z�,�*^?OVK&���"�-�z��2^�tv�s�T"��_��EX!ųmI���wW�c�'�<�.�K-�n�be�e\�
��n���*���B�D�8�q� 4+����q���j;9�5��Q�}�-.���T?b�
��H������E�og��}#A[;̏7p�M4?�1�TC'9�iT��������?ļ,i�U�%.cV�M=�u+.�5l}� =������R�#����"�ۅ�x(�]y���ַr3Aa�K�-����U��RP�wx���J�iquf�q�s����w����8��ʷ��0��s������$�T�utqu� Eq�����*�+	�	�[��X��L�̸<�����C(��-�u�3Rz����P�x\�"�� 8���1�`!�қMW|�D�V(/�]{���Ce��v�:B�����vuu�v�S�%��f�53�KR�l��*��H-�4\����N���	68y�9-�*R-����^�d�����S:_�
Bb�Vu�S^m�GEא��&�O�ʳ�o�䮓p�nhǰ�ϑDڬ��I~�	$�o"B�
�W#��:
͘�;�G%����
K")�E.���Y.��j��*���鐲UE���G��0:GJ�oo݀T�Y�@�Z��xG�����jw��m�'��q�!ɯ"������6y!���P�m���L�xml���Ց �	��Uo^QtS��B�f�<����n3P��^{G˖]9���Sÿ�D�?�U��n8�mp��B�E�SJd3d�P�����y������Q"���|�E!���������9�2��&ϰ�]��/'���bϪ2,t�Z3Q׻�	1͈��i�eF�b���=�=��Ѣm��q��1�}�Tb2����n�z�8�	1+f�?y��i!��,��F���������_�Kȏ��+ �<�s�ֳ^;��Q�0������W�q��'ۜ6D?�i�N���1H���xF��譳^T��W����Fʲ%�m����q�Y;�0t�ܐ)'j����&��l��_9q{����f)K(�1��óȱ�F�!��7i��?����_ԗ��e��{h8`U��F>�I��=�]�2g��I%����
�A�q���D)s|q���ŧڠB!�u�Rn�&�W���7���˿�e���v���G���&;�r\�ag�ūVֹt:E6����C�G��j2��0��,��7X�]z�k�$���$o�@�M-��]čU��`�B1�4<a�3����ڙAa�/7�Ԫ�[p�����p����i{+�1��V�{�Npj���m���,���n����Q(f[Ӟ��O����G�	�ܧ�{�ᜍ��5�BcbPYcR���*-�4R 7�M���Icc�Z�6A'�J�_R#��x�㲨�%��Ն�R���M��H�2��,_�2�+*���?Q���y��4�g��R�� l��Z;����´*Q!@����ٗ�Q��*?��0΅^\S`�$s���Y����Y�k��Z��q�mG��-�%�@�)��#3O��!N��
��YK��ٮ�-�Ȁ��̳�"m���m:�І=B�
t�|���;c'tc�Y'D����Y���{묻L�$sJ6�?�4�
�ŋc��/����}��
0��Ϩ̳����<���j�J����h�
��wq�c�9O�5[�پ~���)�%Z��> �����j��
!��-�b�/��U����K�Bu\��"{�@ds�O`ɣ4�9|�Y�p]6Y@Z���۱��h������sA�[��Fɸ��c!��.���Hҋ�Xs����mh�rX(ŝ�p�Ep�Ύ]L$ױ`
��h��s�k����]\�A�&��&���(�"�&b�֮��F�sW���kD̒V`gڌޞ�t�	�?�v�a���%�B)`YU����������rяq��9+`�w����� X�݁�NAh*�d���Vҭ�i��	��u�q���=i� P����SD���ڤZl jn�6�t*��|
¤��}/�7s�(uM�,��y��cŗ���7uϒ�z�1�mvZD3��xX4�N��\ 5M�Gij!?���q�&(�Dnړ��sa�yV���ʠ��؊YV�`��K��zØ��Df�(� ��H��#:�=�-EZۮp}��M:Ʈۨ�ƭŶ�3����g��#Xc��3���g�c�C"߯�[�IUd��9D���zN�+rh�sc0�p:��5�� �6~)����+2TT��w��k�x��(q|o]�0;̡�),��H��������a�>����b��+�B
Q��D!��B�%�e���x�GF��6m">��m��FE�q(,0��Dw�&��?�/g�/��Х)�^h��!�[z1�����M�K�`�l�RN��83��	W���A��L� NN�ڛ�kƷ���ڕbέ���I��?�51�(v�L��͚����%	T��B���%�<;.N��D�U��բs�l�$��nt�}M>iMl�����D�u���|r+�(���O�!�0@���pq]x�[^�K�������r�:�)���r�݀;io��ĕY]���66q�؊��C�E�N��
b�,�NBR)�I�Ti|L����+�pr��%0�����U��v.�0}�[9�aY�6�5k�����vH�x�(R5�3F)1�Q��<��,4Q�}���Q�jՔ��"-�����X�y�b�Q�Zy(g��X�R)Ph4��_����C�4�# 2���S�j8�� P��Mz�\�Oh���(�x��D�eeK�22��:�	�%.Z(�о�[[�S0� �)�[�ȗ`�LH��3(�V����"J!L�v��2TN�᢬e��<���[
>&�9B�e25����a_Ts�#]�b}B�I`�j���Nf�1���֛�p\��,b�,g�����ַREL&���d�'=e��F���]{��Wf����{����$�*	<���7*^���F|��	���7��}�fF:�ev�c+@�=L@�L��k�ie�p+�cZ�Ϻ�js���cN39��	����yC>� Ը³��(Ҍ�y����ԑ�]�5��銵$H=���p�pmm:\:�L��~�5Zl�{�A��r�Hy�ggwZ�C��R*���ތI��[LW�x�2TZ�dֿ\}e;§�X,�WjQׄ_��J�a�]pŴ�.�x�O��V�0݈P��މ�-�������<|�gH0���j�.�8��ǇJ� ���۫*ȉ�ĸbgp����I�k�[�W���}p8y�#3��4�=2QY�����oyw�>�'Qi��(�>t�T'F��ş��9��ǩʤ�����b�S�n�0��NW�?�����)cvĎ�m����_��Ge㍂RK�3{��E�w�S��u�����dF�d7�]�!m�s���n����.7���')��q z~&�*����f�[�_�[��f���� �!���$���������m�M�2�SJ���S~a�\^�wE�����*�� y�����LM��/�K�l��M:����.�0��Rҳ_���Tη���;�}؝�o�-�R�}X�7�U�I�F�&_=��Ը׉� �H�Y���=�:�K��Wx�y��tn�*�ƒ�Z�o�>vLM/����g;P�����֮���^=��'����La�r^�����wk�r�@���B1bz�e��]w ���]�?P���3���]�b��=�B$�� ͂�������'&�y�J� X)���N�t>�	�ɮ��n@++5N��S��G�Z;��ސ��Է�7��2�����ܢ��/��y�[�/a�<�_w�-��o�;�s��m�۞:���i��yCl?���A*�U�C��0�}�|����~��eai$����rU�/A��9 �8�r�²l6��_FDt�$�>b�T��?z!��H��ҳ��~Uh�P>��y I8/A{�n!�qY�Y�%m��MTͱ�ޅe���J{���0[���k��k��g���_8mN���m�z�P^�սҍ҂���q}��S.o+�Ɇ@�ef䅎	@�~AS��)JtC��S/[����)J"�V�������Rrs�ӂ�RZFʨM�r�k��N������[b�*�ͱ��5�i��Z�:�����}��)Ns�!�v��!�r�/��e��������ꉈ�'3�S`$���l���|x�Y�$�TS�6�!Hc�INh.jv��K4��s
�"�oh#=���Q*Q����|?L�8si��yL$���$>��s��O�\gS&�d�^�v����мv�~Y��� �n+�`4�������w
���MNU7 ��1�j�/�(����
-��R��$�
tL7�\�;�l�ZՁ�#h��
䵖�x$[�7:Bь�l�IЕ���#1t��.05�;b/
�% NP])Ѕ���'�V��T`<x���\�{xJ�%Q^�e�z)�� ���x�*Ji�c���E#Ւ-��l�j�����Ƈ'�rl�_�3�	��[�r��-������ƣ����[�M�"z�8]"�!�k� �נ8*���#�xĵ���k�����E����9X$���W�/g2"���^b�@�1�M�ٷh< �����Q�).# 껆��ɼk�c�[����F���r��s*����E3�]$Y���f�GK��ӎ�of���T�
l?Q�u��ѼK
���P6���Q{���h����4O��pi��/� �ekz �6��qio�����5~����;����*��Pox��u���������8c>����;�)r�0���>O)��B�����>��U���ߠ(YK2�a�����H �O٪�7�_m��_܊"ܲ�n���=�3�b���;>���4FE��g���^}��q�O�I$�q�Tn��tB�--Le�m������݉Z�o7Ȓ�鹁�F����	���d�iU�e�)�^� �
A��������,�4�&�#�A�����I �wKۨy�N�6X�Ybk�K�k"�y�0���d�"a�_������V~�k��!*�}� ;)UD�镌���b�
�)��U׳A���6�҉CC٦(Gm�"!y��8�%��
�`Wo��*���Y�N���ұE:aۑF����@�� �+(�x�1��N�*'�Dc`B!{h}���9_�h��
e��P&Tt�6��(�ʰ�f%E�űO�g�e�)�;�=Z�;4Oyh��1�-�x��V�P�z�1��r(�@���xyM�v�R�n��h��R��ܬԮtt��������8{S��a*�X�N���Q��-�&�	�����fd,�4G���@�>^]�a�\��)V%5�|x����������#��wa~��6�V�~nE�Yjev-7��e1��e(��0V��6�^�����	�H�x)�Ie8�[�RI�����o�G�}M�W=����6��]��`8����
_��3��
Ddͫڰ�A�{G��'�U��G�@.0���#�v>i��W���\�o|��Vg!��'��ȁІ19]\#O`�6�^���LHb(n���u� !�D�ؘqܣ��nV"u��=B�$�\���T���;
X��P.$Ÿ',��! 
�ifL�>np����0�{��������>J�f�?/���� R��U$3\"Z�6��SU�:��f�U���9������ϢW��GyP&�\�@ׇ��IT�o�ӌ=u�8Of]лЎX���s!h����M�"�_:�z���5�AHջ4��!ݼ���"}?RwBCD�{'��^0�����.,fɢ��ߚ�Gr�����p1N�Y�	@U�F�i)���HP[���U7�F8���{Z�˛.1��!+����*�p���rҳ�;�&���"U90+IyLcNvKɓ
�y6-�)#B?��a����B�E���Twُ�$����[:�w�̃o��X"����V�v�����5}˴���������S���VR��L�a�(ōK;|h���/DօB��*X8�{r�U}�qli	��C�t����;,���Ԕd|r��k�#,�!�܌����or 4(��Q>7�BUl^�p]�m�~�{p�F��%�D�NPC�tĪ�#4�'�7KR�. b^��N������ �Y��/=�+˹�c�Z!W���H�4�$�8���U����+[����ګv@��w��8xkG���� ~s����ۡ��̸�m�Ѓh���*`P��b��еL�ZV�`��	�0QQ��v<�Q˱�x~J��4�[r�peU�s] aE��\O`#m{�@�ێ��^�i
�qv�*�MU/�1񆋦)����y�Q�N���d��n�� ���	�AKٞ�.Ԗoz8b��2=��NAab�����o)E\ŉ�X���R����FC,T�� �*� �q,.�Y _ �F��(��B�L.D�%7͑�9��L�D�+��q�S��8@N�yB��o�qƪI?n&B)�,��TV<��Ug�9�G�����n�v�Y�d	�;i��3+;?ߧ|����m�.��s4�p����<��!9�((_D�i��W��]Mφ�����.�Y�l�FHR���*���y�-*k\�\VC�֦�S����!�b�<���r��d��$I���EI�K'�����U.�[�v�Qv{
A~I��5�}�e�m��Y� @K���`.=~#���D#�{l�.�ɯ�h������Ζ�飤ﯟ�-�ʅ�z���g׃C�ZV�Ѳ;�k��-EJ.�-�3N�3%_�����>�Oc�?�53Dʗ8ʒ���zռPt��e�,�F��A
��Y�Zj�n�upޏ�v�]�\tV��@&�z��Ȍ
��^Xu.�7����E,``�>�����xI�s�K���[?+=�[�<���nb%�)\w2��_��E��U�	�H=���c�i~ӷ�Y&u0��)�K�kE�����U��ĩ<V�7��K����q-����Ά��*�\ڐ��� UiYx@2y)_g�
t��n�H\{�BX"��8�u�^d��kw��(VH>0��� rЂ'�'&�7��P��D1�U]wX�9xm7?��9�����R����@�
��p����-]ɨ@�w���������{=>�M85��/���ԛ(S��Uz9��vV���n(k�/���X�L�ql�];��L`�"��� G ���h�lA0�҈o����N[^	r�!}!)5�H����$J��Dtz�����E���`�~���F}��Q�T���ծʓt���� ��>��T
���Ѿ�T}0B5�0Q�#_C���}�/�P��8�����'S��&��-l,�Ed�U&UM$��jvw0I8�m���'S�	��]���8ɍ�t��w
�뭌�}2�����h"��.���R�*D����8V���I�XXCV �˂{�����^a'�<"o�^��\�Q�ׁ|X�3(J�� 	�o�����=1��Z�toؗ��X����0S�p���{&�.(� s@"�3�T� Z��׻$���+յp��E(5"��X#GE��LP�!���(d�'Z��=íp�<*2AC���)b�����ncd�N��}&�zWːv��o�o��F;0d��$���	'��Ղ��{��	�np,�i�C-F3ؼ�0z\/fE�t{ܞ��V����\�����֨��w`ȰI���	q7����<\dP?�f,^�`R�-�\Ah^�ڈ�(Ф"~9�?�1t���0U�7U������P�<�2�Ք٤��5l�1�_�@�%Cj����͗Lr��� ��Q�cM���;�QI��PRZ؟s��0m�8M [uq[%�<^*���l��Ci��%q�oJtF��g�.�1}�@�͞=xT�ᓒ�W���?��Q�%0��o(R/�$ԃ�&uV;��+'[��o�������y��+��-`.ğ�0���D/R9,fd�s=`�9������.J��V�`�)"�Q|����4�G3`*���jʓ�+�U]�,������T/�Q��"�3�rM��<,yڠ���2%>�E��DI�ፚ��Fl7�z=چE���[RU1c�]?ّ;�(B�{����|��vT���#C��x}G=W���I�U_d�e�h���?��فD@OV��C��,p������6���4�����#����!BX��P6 �XzX'���}O^)���ˠN)����A�[��$�65>�u���(@Rl
�
-���;T����A�XhQ�2+"��v��
���M��j�5���%��ph�����{�*'#�R���~�2����-!�F����P~���Zi���1��-)�_gJ-Q,�9Ԓ���V�m��}sLҴ

A��:�5Jr�\�2�_fD%�Ons&5�w�;��f�����P�h�>��_T3	���	�D@�������^��>'��՟�?H�~Y���f��=iC����t�����m�ɵ�q��oJS�E#qxG�X%H+;�s�]c����Nq[G&���|9��h�k�U��@�l���]�7\�9�lݖ
��qc�T�}�O�� <m��4�6�z�`�_��
4�MlòhM5����0C�X��B���!|?$d��>Q�z����e�,A3J$��`7�w�d����~=;�,�B@�~���I���{P�`�����$�1�����Ц%�@gU�����\DzRo��#�I�6�ܡ@�_r�Ȧ!f�XiE����Iq}��V�*��1��u���O��б���`���Uۯ�8��,�N.<"1I/6�S�u���������C��`R�
��O�,<�o��U:֢�q�Z���@#�4�s�hr�� �s��`h@i����N������ڇ[K�6��$ۭ��J�=���5���*�de맅�>k�}c4ֽ ���Ͼkf������	$X���"��]4־|�܇�
i�xF-��%W������3.�M[T�@オ�K�+X}[U�C��L.�8�j����Vνp�wB-���;������hT�8YP�k��7�4lv���'m��6=�	��V�mu���#�� �R�\�R+Ȗ�(7�s��oDy�]��͌�Ն���P>��63��i�8��y.�Ӎ����1*�#����en���^".�^��1���S�Ah�"����J].'��˗t˫鎒E��R�%������{��x��cb���ַ4��2�^o���-{��!k�A�%ooN���"Vr�����?,j_�:1�~�Z;|�ծ\���'�N`���v�b�R��
V8�[W��OC�#���ǯDc��mQd�k����a�r�	Z�������]�nEP��^?��<������:�j;ߧί���m-��&6@�Y�X�Q1�z[���;�P����g4�Z�S��'��4H?�R�a!1��3N߳Y��$k����Em[	J�nci�����c��]��P��_�C%[�f�%h��y��Ty�N#�;��H�a`���~�'�$���/˱>�h�)�F��¶��J��q���H��$ڠPmO·\�[�V���=z�#�b�.�1�Ԋ. ;��A'tZ�TJP�f�+@��C���
DQS_|���9��]`��|��O��G7��#&^��H��<c"Ue�B��5%��*ExRX3�@�A�i~��O��Z�v��X�(���W&1�}Yə���
# p1�I����q����dξ\�lFS��(*��.�$6]4�G�ϖ�D:����9Г�SƄ�Zg�H$%p�$���A�c�f����%��)�eKV����7��DXu�99pv٥`����tJ�.����:��9�{�D����T�������ڱ��bg�t���f+х�&2كe�P��Gp�C����*=��x��n���r*��|'��,oe�V�7���	2z\��0n#%�a��2կX!�?��%�Mt����>���������e�������IxPT�h'��x	YԸ����
﫢�bK��Jst��X=��1`y�5�}�ͩ@�)wL�����%�a�J��Y���i�9���`�P��K!�o9Mr��wm)����6���{�:�$�˳�<�d�6������i�8R�.��ph[�E�����3���0��@��ǗQ�ӗ7������P���G����7M0�m1�X�E��.�S��]�'�~�ŀA�x�����쿖e�<V�f�85�_��&��0܎. M���e�_(!��x���p��܃?���2�&����P�J�����	�X}5��:F7b��C��j3+�:�2@��w�Ѣ����D�rd�-"�C;����2k��
��jnv���|�V�O\qCY:QtF^� *����C�{���F�|>�~D����fH^�ޜgQ����������Ï�)�f+��bd�⻂��?��.d/@ Ry�}Dv%Z:��܄�`�:^H�h���6�� �u�M����	�O�'���/PBF?�*i=Dۃ��r�ɝbY�M��!k��:ƻ1��Ѫ:�OI�^����(���	�]��TYV�ܷ�C4�e�1�+�P��k�}< �M*���	1H�$ZuwsKC���9>ޓ(��ԩ@\����0rn͆hb�L�S�������c���[Z�k�1�X`��ߦ,QR6|��g���d���?���N��y+{�&'㽍G$�聬�������o<��Ǿe��l���b/R�{��.!��0@���:���i�|��F�-M�_�����E`؎Vpa�..q�kq{N�,EO�"�y�����?ּR�J���L�*	�l
 ��d�&�����~{�z�KS)8\�9%"���;��D/vS�y�l���-�y؛�j���S2�W6Rߵ@dx�Ή�5��b�I>�bG�y!�ѫ�.��j�s��rksҧ�E��[�����[`(RR�*�@�F�<@��G"�a�ވ+� �y���j��}Z�l��ۜ�`����Gtn#M~�ʖ_Б�R8gi�O$��L�	=��i��K=����Rx��|<�C�;�H��!q�{,{4��"� ���g(գu�!MX6ԋ��S��k9W\+�Pʊk�a��X�YW׌S�
��w/�z�h����8�������a�K���>��W� �C�@6�<Z7���������-�@7��,PAF�S�"��Q�8��J�����ү�-�s+,�!�����
_���n&]��z9�Ko�y<�-QUK#�Rr�Iq9��Zq��3�N� ���h[g 3EJЯ�E�O���2`Ɇ;�]�T֎%ŵ���������)k��p�_P���$�m�v3�2��+������'�D�G��`OUH�XL<�@ZL(��q�-�q[�ub�|�NzK2*'0�1��P���'-��|��}Y2�?\ rU:��Dl�2|�+�#^^����%�
�ٹ�c���\���b��DBr�;�#;:igV�����4�x���eX� YR��_��u����w@�%��厠/�U�Z�H4\F���`/���`.�;M��;P<�[ �,lm���g� Ȉ�(�̩a��3Ҟ5.�-�Ⱥ����5m�6���'���Dٌ��Y�#�du�1z�Yl����8��+f�'Y��9�<�>x�Gt1�~�_K�(�l�u��5�K�����\�|r>�ˆ�*�gy-/S�_u�yN{'=c �0��"�i��5��W��y��k�^=x���I�Q�,���������I 9�r���-l�F�|%gd�~�9x�\R���l7��;���+� ���mzN�e&���K����5N�*n5�Y�u�����_��-�K)�?%�R���^�������U�݊�TC���/���)/�k�0ʮFk�]<��2d'q)�[��`�ÚbYZ�a��������TA��3��u�cY���� �A�T�?�� *�qP<��,U*!H_����.�f��/±�/�yI_�fH�g7��k�!m�9�뾑$�Q5���N#������c����B�_��t��^Ͻ��3�}
6�V�T^�����t�4��g��/	<b}Թ��gwUl4��I'~E���+D��q�
B��#,�����v��Ē������J��Z��I�W:�n.sw6��m�����~�]=�*��r�1����@ޱ[��1��D�D�A&a>�x��Z9q�D�n/�V*��@��p��G+%�cSv�_�����B��\�x{�23ÓjMx��zB��P�o�P���0��%�l��Lr2�hc�������%�m SK�@���m�-p���K�$/<q��M���X=�����-ݢ�~���Z���ڸ^kK�F��`I�.1
Ѥ�x�w�/���
1�Z2��|}�?9�Y"�����`sx�9�M����f�]?�x�l�6ՁTl� �!��@���4r�J�gψ�l�x]q&����R�h�g�g����|53��$!�2��њ'9�>ĳW�ˎ鰂���@�BP�5Ѵ�+�9�j��W7�Ũ�<��odL������������DC��{�ѻ�އyV�K%��>-ZIl�%�������Rɿ�1�R�  H)[5m��h�NH��ג�fĺ?�ѩ5�L��\��i`�3��Gm�z
��r"Q�w�̄9P�Vx�.'��]꺫\�������U�����?��u�VC7�Te��������I�����v|⦃�.�_��Kb�Q�����8h>q T����R272%�İ�4PtQ�qVz�Ľ��E�A���Jɢf�`W.u4�At1�.��؅��X3>�3�U�TY�M4�C�Ѳv}6wdW�:�˓6�"�'�e�yB��P<��á3��Ԧ����Į���d]fLwւ"Й�bS�<2�ԡR34)����6��R�*GYy�Q��Jv���x��YR�Z��y��47��[����A4F��͌�@'�ļ�0h���K"K\�M��i_��Z2�G���
7�aiw�g�~NM��~�`��0��O��np[���{�;S��Ǳ
���g���Yv��KȨi?d����`~����E�)�A����E��5�f�6�<��W{�D$����xX��b�Df��!��K��GCM��aY�O���� ��e3(D�˦^�\1�Q+��
\��Tᵊ�]J�����7O�_��7 y�ϭM��:�]��������������µ%�'
��4��R�M��	=�2u]F#.��q-Y��*��� ��Q�u����.}���]��ض.�ʀS����Б�BzA�ӡ4�3d%9X�U{��fZ�U�:���J����+M�'�J�����4��v�v�f�"�
d$��.ػ�o�
�k9�ϏGASn����1�-TZ�	�:O}�M�l�y:g��!Q�iߌf����^�Q�6�3�,�ʔ��(ִ�ہYA��;�^hS���a�C��O3�R��w�CAO�Y��Bq�i+a�ؽ��z&�
#Y,�v�a2����seGUgA+�If�����5��9`(â����q�RV^yL��;eEp��ʃ��9]y0.]���쩲K��a�D�p�[5D3���1Y8���S��ѵW�m���}��.���t^[F�Qe�kI��!�;"�Ӫ��n��1b(%�h�so�w�?]ʒyn��I)��k��*��t��E~
�F�C�G�F����T5Y�;�(=�Z�'%��Vp��V3�Zƚ|?�f_%";Nzۂ|Vs9*,
E�(��rE�>�v��%M]�Bz�/-�N��~4+��=�Y�l��H����3���`���*Qc�~ScVI� K`;X~S��*������m��9�{��ޣ����]gls�=�C����0#-{I))�3��%avʎY⾚��\��1��Ԕ��f���4�֘_qE����4�Z+[�ӻ68n<��*h���!^
�т=��u�O�Bmj����=	��>�W6O�֎5@�tEZ�3a�C�k�I�ʥ��3���4���kO� �}҈�}��Z�C�o��LwC�QQ$g��1��5�T������@����P�`Mi(^���*����&�whG!�r�ș���u)Ӻ���?������gVb�[l ���{2��,|�+l��Gn@�m0H�-��D�N����D�@K~�L!3/= ;yt�-�P$���V6�֨V��R�/Y��^T�3�L��fUMx��\W����:w�yK!헺��:~$
�E8�&�.�Eٴ���M�c�M��$*V��h-3f�بi6~��m�udK���[��\��hǰ�C;�D�2yT�~��&��f�2�0a�U,�����1��8���rd�B�%h	uB`����1�������=�9����f����N>~�e�B���H<�q����p|�Iy�SS�����*��\��}��
��:��0�N;�p����~�کpZ��u��[����HCdu�)|<H���{Ė�Į����q_~u�B��{��X�g��cm�|�H|�4�K�|�6� �
�l8� d�}� &G�孌ziߴL�S ��cx�I�B�C��r�	����žt�x�8�xʓ���!��;�F@��3$2z�t�$���
E�M�����PePq �U�Q��$��<TJ��i�x����J�d0���B�/�����VbЈKN�x��y��z�K��C���]NJ/���L
�;l�H،�����nÊ~#�T7W}����	%�#a�*@RM�U��05��wA8��9��D�N�f�nv�[vAd���.`�/
U���_��Z���7�h����j3��p�y�	;�U���JhV�ߚ��\6�V4X�/|���"8�uπ�ے�qXu��郎�ދC��%��X�6΢�(����'��Z��?
��T�^D8ԒЋ����~t�u�u�f�4z��E��3��D1�H��T�j���e�R�N.K�����K,	E^�S?�a%����Җ�6��n���}[�V<3�9 7n��N������q����`��0k�B��=Mi�)4�#�ض:nu���yҮ2� � om,�aQ2��Ӊ�<�MR~y��(Z.��QԼ��)e�{���l�!w�䠅���d�aF�%1C%��5G�`]�>�y[�e�������4��bc�׆��V	�i,Dӈ�JP��^`3Or�y��;_��Iq�8���㢓���L�X�����)S��^�C��5J�JQXCU,��Ԙ0��$k���P����h�O��w����h��?L�8��<c}��.��?+��{��ڮ!�����j�R���7a(-����6p%��s��s��d����,�$��m�np��ݼ����Z�1��3��>k>/�,����L�X�����\�
��2�aS@� �A�)w�	�і�x9��1�`��42Wr�?�-�T���u]c��پ�����=�v��m/�� �ͨ5����-�<`�:�@�4᱾��g�B��0O��2��Ri�&~O%f�I4���g��M��>��X�r��ўr~(R���K,���80�G��sJiC$)���P��'Q�K6�$�z���%�(V�f�KtG���R@�y+�/(����«�6�vǿ줞�@7�|2�|���:�"׌��WB>�(D�ʐa���m}*��w+����M���?��o4lD"A�T�X�.���c���ۼ`�{NT��\]f��� �.B3�<^�\�H!�A��&lIj艊:�=NT{en�9�`���:6�M�+fp��#(Sd���Ѣߤ+X˚�`�ԫk��p�U,C#���������1t��TW�Vς���V���'+�[��^�y�Ŕ����atJ�����ޝE�5`�
�8 �Z��,;��Vz�D!��y�k+�:d��b�M)�uɽ�W �5��ݲ��:�)r���`�N.�2YFb�B�@�e��<��pTf�ocO�@�ޕ�.6�,p���⵲�*��¤7S)�Wŉ��:�(�\�@et��E�󎵉'�,산�c�6�b��Q��|]CcI���&ʒ��X��>��i:p�w���J%�G>��y�R ŋ�
�d�h�1�,'q���-��&���X`gR��9R���?R��2�v��?�V��1ԏ�[�ӳ�@��% �gUE�|��q�䊄�1q:"��"��Φ���Mba���վ���S�������Lx��~����D��#-I�� �9Z��>����xXw��� V��t߁�NGtH"^���Q�Ł��mK������a��ꤕ��Z�I.k��n*O�$C�
�¸��$�$��U�úL{��f_�>���=��5i�����'<:�O�	�ZϘܨ�	�ix��ںCu���'	�n�t��H�'��gx�?ΊI�gu�6M���>�U�&��崛���*�q���Xe%I'�3���I9�a�O �BՐ�V�^�B���9O�G|�(��CT��p�T�FԌ�>�9Y��|����I�*�d��P������;�ƕ���.B�M�A�x'+=t�4���ǐ���x�̵l��,��@s��6�/�T��1�5�ϸ&�>�oP_��OqzU�'s��jW�O�u��~ssK�n�q�23�(�[Y��0���1�5��:MK�Q_A+���u?|{���[b����u�2����'/Et�m�}`E�LX����PzUpj�^�̠6�+Ex�϶�BǑov4F�^�y�a p�I3�����<�_MC9,�8�JLm�!��1��X�>�V^�Z��DF�9�~�p>��`\��ڈ�.O'���������CWA���X*C�zl}�hap%���G�OQ���2Ht��abR���oZ���ĽR�źQX�Hz��ȇ6J��Z�WW��¯;5�/�vgp��K�@�j&�o���=���ߑ��c�'r�5~#�PZ�{2�&$�A��gW��Ɋ�,������Kq�
l�h���n͋6R�6éY�vG/00X5��@�Jb����`�NH�$�SO�W�v��ɮO%�qY������EZ�L�Hs� `@XͿ�%����/�7�ۛȄIEDm�=ˏ���H�o��!�k����ABa��Zak�f�֗�h�������8��4��o�oܲ@�.do���^X�[�YNY`B
:(j���w�_	7n�^�V�Jɜ1�&���í���]�s��+5ӝ��^�j���~�oA�iک��"�,&�C��:��ׅ�Y�VXf�ۯYn֯�2�>=<�aT�.^C���n�}�n��ċ��Y��"�qg�=(�d�$.ż�>9ڝ�&�?��`�bb��� H��t�a�u�`�{ZY�˻�l۔b�w:
v�!������K��Hb>���9k�������ƪ���+����ZV��6I�%�Y�x��S� [���i��Y	�����郤�M�%��e[@	>���j���ZzDlI�C>
G߄��]�M_�Oo��5= ��d�����=�X�;e�q�X��7;�PX�\z�l<����\��K�}������F
�H'r
΄����S��aQ2�r�����f�F7���t���6����&��*P �hw�}S�����ہ�3�����w�˅x����%�v�jL/�[
���Kj�:^c*�҂��Bp�&����4e��e��gⰓu�]NY�oC�ȟ&��&��eM����Q�0�S��&�^��6+d���,b'z�G����N����}�{嬟mo�%\���KJ����͸��/Cv�:C�=+�'i|gمT�;]�[/��t2M��;�G��K�E�|;?�R�k�_7��e�V������
���!��Ӻ��ĺcg��7���!H�}���-�#��(�I���a�zs��;�4q�	Y��};�G2AtF~t��|=�M4�%ѠE�KKO&B8��>a�s�ө[h�����R:S�p�+���������CMߠ�KХ�"�L���V{����P�s�g} ��F ����A�g�>0z�K��*��.!��e�]�X�Cޢ�M��@���^LR�=Y���S܄X'�z摰u�k!�@�E�#�eL�~s�c����L�#&&���-��G��Se�?�D�Ϡ$Md�Q�S�{���od�[�\u���J�u%���^e���ʘS��h�t���-�Ld�0M�Ҋk�6X�n�җM�9�	p����E�t=W�d�В�誺7��B��se�8��l��Gʶ/$f��?���1�0t)���ZX4���Ŝ��L&0�$�}���s���g$���QɞI�� �ͳp�M.'�c���B�mL�iVJ�H鶎
!c�kY�U��B���U�%.���l�q�ǘ8�VxƟ�3�����E�����qm8�=3�N3-�壻_؄W$���Q)W�9ՙ�������)B�F��/��YN�Ky�]�>2Z�u:���|U��r�|G ��,�h0�܅+z����
��Y�60*�hۖ���̝�i�#O|�ߙ����
�.#5�I�uNx_����b�I�c$�U~6�ºTѧӨb��g�������w��YZ��x��mNi
��-�S_������Ȗ�e?�ȇy?n�&�e� atq,��Y๜�v��'���v�n�)>M�3���s�\#\�Ͼ�F+�T%р�`Å���6�������$LI��oՒyI7wf�����+Q��"X�c���Z_g�z8�(�-:��`%�7p:��b��%E9�EI�Y��%�<�ɫ���� �@��(��G�}H��ރ�R�Z\�>�M9�!��z��]�KE�|EL�R^�mܪ@��'���ʓ�	��/�+�oMT.�y2L{�������R֯��t�ÅG	��;[�*����p=�	&1:.
o튶�Y����A!g~�me�7���'��KH�r��qa-Z��oBI�c*0�h���5��m]s�Α�ǿ�X����B�%����kF����>j:���y-H���P�4)�����?9�v��\
׾9T��oۧ��f��j�1���]C='�s���ݝlb7�o� J���[!J���}vQԈ�xkr��YR�]	n��L �)A< �Ҕ��2 ��٘�A���		��ܼG���V�y�?���S�~}��CgDŃ�����.�M>�bm8L�0Vp(������x���Rn��4�h���0��ek�����E�%q���Ky�|(��0�k"bbu�v�-�U����G��4��k=��s`.�)�H��oPaL������[O"�������UYN�P�c�*�'V'�)����-R��y��ٻ�����QQUhKb֝�c(H�'�k�+�1T��i"߲�% �ޕg�rf+�wh*A�+�(x���C��rs:�������z9
�ASf�Bw<Wr��"=�09�JS!v�ʲ�s��_^����#4��)� �W��<�G�!�(o�<~�ZGׁFd@FԂ%�J}Ʃ��fm62�h�� B_&?w_�ڄ��'qE���[j/X��fo�h�� ��K�:ܻ�F��F�JZ�|h��
E&�i;��Ћ�B����=�S־�����|���j���ȓ�+��@�O�4�}(���s��N��E��c�%4ĈӔ~����Ў�;�ZXe5=���mDrq��U�v0�-�_q��lH�ٲ�� �}G΁e[f+�������֥3���r���֢{�8 s�<��9r��3(���hxi\;�l�p8P�蔞��Lw5۷�͉����B���w$ַ/�9)��5��e{R{�sPSʷǣ6�S���"U�B�#|!)�-Nܓ�i
1�n���&�k�`�6�k�f�k \똦��&s�Aw?(Nl�bet����T�i�x/�*�3"꣖��k���hđ6� o��S��LV�ٸL���;������t�+6Xr|mHw�EK���I?�CO�n���m���G��4F���FtEOLI���ni[۫�aL#����_%�V�Ch$�̪�1ak��"Ǐ�����8k0�ڿp�Ζ�ٮ���`���;'�萦�t���I\u�t㸍T�u�>be�5V�ae�]�;n+8uJ�I�W�CS�ݪ��0�5iz�BgE�J�tb�.�n
�e��)tl�k�v�����d$TbC�+s�~��4 yLXI�#*�!�KĠ/~�~�֟�X���nX���&ϫn"Y�aF�����o�o�bE�*����L*���y�v�݃�� T�VVvM�}+����
�s�����a��r��p�T�jb�4��YR����H��Ara6I��f8Oڐ�fJHخlW�C�_ڔ�o�ja[��+e#VI���dޘ'8��E �;���
&Y5�˯�Q����w�+ ���7��j�`�����Ŝ�dh��_��H8,X.����ތۑ㍼�jE@ݰM,{[r�*j>���xB(���BjխP>�Y�i�u*�ɟ��Z��)ɼI�[�D�+��4,��~����c��$3b��$Ѳsh񐻫!u2L#��I��t�� zg��#u�Y�J1H����A�
�#�pdI:��03�8Xk��5L0L�rs~��mÈ.<l*l������,�D5߹�������٬���6sj���R��6�lƜ�	UB�t��kL�J�r
p�)+��vw� Lq��.�d���P�t5Y����_6=�٥��x�x�8��hqA���&�
��yF���t�?6.��W�z�JB��2�iN�(���a#���-聸9�Ӄ��	a� ���m��w����v�$\�����ߠ#�2�y�?���z��lBvd�����·�n�H�ɒ��bᡓ>�����w'�*ẫ�2kp~��U�ֻ2ϖt�_��כv�9��5iv��m�5�a�޹sV4?Jx�HU�rf�m��Qa�a* Q��Y��I� ����v0��zL���5���t����B#N-D�<�e�{����4�L��s�� r��1�B��7�|��(�aw��*����o�
Go݁╋S�D_0����qS��wl�(�D�x�l5���$�y���um��n<U��BI���B#�l���waG�/B�E~F��6T�#��"�p�;�b��v��I��bj�ҹ�&��������_��@L�$V�Ο���g�ـr�\��6��X6��{�@K|��w���_:��}!�ʷ}_ց��NG~v��r*3�.���b ��e�
L�r��a����-�|�siO�Jzcd��$'��ї7%T�>	�fL����ca�	1
	���1���o��|Ycq�.������7�K{�$���E�r�F��?�u7��&""�6��ͩ)��=Y5�p�ً=C��r(Z��,bZ�K��zV�Q]�p��qit=]/��b�0�f	��<�*0ͥ�cn�x�{�,����8���?�4��L3GSHg����R�?��X+K��d���e�%|�ތh/�7�Hb����Ʒ�t(�����\�_�4��o�|½���T��7Ŷiۋ��R��A�ȓ]"��m&�e�m�/�5�J�b�o��1���y��8�a�o9\P�E�Ф�U_�g���z3�'pbVi����n�5B�2gq��'���e� ��)�Q�/m����a�ʣ?#/��6�g�a�s��x��«�h�ϸ/|!��7S5C�j� ���S���;�b�_J��@���#�p�&�B�?r��e�9����>�ݎϯ�wWv�G�8#�df|��S�^�b"�6-�P�L�S�����&`����U�c��=5J<]S>Q��7E��WU%�ɉ-ě]L�E�#�{�K�F/�)�-.�*�H�&ɷWmj�h�,����z�F��kE#v�m��#��Use��F[�IM�M"a]b}W�	���hn���UYm��*e�����t-��N3��2����P�F��t�����K�N~����Y���q#���0(VV�!?�|�veK�>�l������=�R�1'ͥ��pA�d1
�|*;il�ɶ!���)���2$-c��n��"����-iD�����\H���uЧ��S���{��+
�{(�v31�H)���J"(��V�P�h�G�ǤJ-�U���Sd;��~A�YT�%�	�-2A[("?����~�m�Cs���˝-�Ã߬���~���h���1�s���J���/���p���v�_ihI�(��m�eL���W�|Rxp��K��OE:��/�0�R�z���҉	,��$^�aн��K+=9�5B���d�A\}�K?�{!'����ڤϜ!ia��KPx"�c���uE�?��8�n��\�����y�!PG$�S�i��+���r����􀮒���f��K���) +<4�7��.hoda�o�^�XY�i䥞\7	Z�2�+|ֵ�ۄ� FGpC���j��HT����r��-�I��%J�3���o|�\�sO�rk���)�]���@�>�� |�2�o-�S�[���-"9 �=;�mwd�N�Y����:'$f1��jk����*�Ɏ�7��]�X�,����j>����Cʴ �9�
r������'�q�?z��?��UWw�A��F枴�3֝4,A���lȇ��2�9��0~�?�$����~�X��֬e�רU���(�'-��}� pBN�7�K[�P;���0w�iP�� ��
W�A�7)r��C���U4��0�1ȲD�&�{4���2��� ���6!�bG��1t�z��d������i���\4R�c$��q���\K@i���:�#)ޯO�����pϟ��22Յ���W�e���cߚ!���D�5��e���������?�ѹ&3N)�ru�5��䓝�� ��,�O;>��)�(�hP��ٛ6Q�yNw�������57���3�����Ob2�\�v�]A�Ys_3+�� 6Z�hǍ���m앙6�!��X!��bW����T���%���!4M��RS?���36'�@E�z�����"F+�Jc�r�HS����i�>q��W���<��3������W����rbz�;%����/���T��D��5-Jr���Q��<�Ƭ�p�6�0y��3����3{267�����`K�/�q�1SM��{$�<�L�>�M�,�KG�L��o9��S.X��'�$��m���7�͋�Ux���#)N剨��4��g?,���v��a�b$3 �=2�vH��j�@�9�^�0���(?�JJ%%X�LY~�B�[OA�dgh���Vsg�`�r���^�o4��Utr�/�?��j@�8�<�3�2����r׀ck�q��8$f��%*Rk�g�gmn����Λ�2�]����~��f��'矍z���X����@u�;ql93CXKf~�m�ص��/��a0-DR:����ۘ�����]5����k-���cD��?һ�ќ���w���[ 얬�@�<\����w9��3�_:F�nYb�.8R��j��SH��" .ZP5f�+E8���)�X�{0y5�Tpٞ���c�������2-\��S[ܜx�Ҡ�xS_"p�v��o�W�I4�xč^��!�� �Py�6Cڙ�ԣ�̤ޘ��7���r��kH���[�f@(!��^���-Uz����8�|�t�@��3"��"�Pi��v"��IoL!g����;`k�uv�V��J��Qc���+�n�06�E:ͯ=�V-�����zZ�v6�ט��&���۶:���)�z-��]�5�w�J���x�T��3c?c�U`����r������mr��mڸ��?��~"�I�w
�c�Q�r����A7ϴ8��R/DE���M�1?7tD�����0�O��B�cnq\mI.��d[��$|g�=��jl�s�6V�Z쇳��6>�����_��N��;���/y��)z#)��Si�z��g~Zr-{�t�k����I�+�ROe#�ӼE�d�a�����d�)���1�l_.�H>+��=y}/�%��}�(� >�JD�iU8=`��hPr��@Q5إAN�r&�E����.'�o�^.�<�^�H���v��Ђ��U�7{j��/�����WE��E^��������I� L� QQ��^���/����
�V	z��n��]�.u���,���t�)k�Er�P�������B��)R|�(�{��&7'��"�Y��|���y`C�7�ѻ�! 蒋$]���޾���0��^�ro�'گ|�}蒟u�6��Ĭ�7�;~�@�f��Pډtf�C��qy�ܩ�|�ڝ���1()��	z��5�ԙ��J#��V���u���#���,��d��[y�4�N����H����)�x���v�$tתݕ7ʞ��{���kT��۞���K���Ǔ;P�����'7Ֆ�?��#�o�T�m�Rߚn�F�9_l ����,�;�e�=ݲ����� �����	�L%��+m�M�70��w�a0�D��{�00���Lt�qA�hwg!�\��C��Z��B���F9b1�spD��,�����d�0��C��VO2��	K)�L_#˭ړ;�����)��d��kn0�){;a
��	a�\޴����e��
��_�h{�/e`rSF�|�	\�@��߰a�[a�;�r	��Ό�I��|T�*�X��e�WI�5��I�G����,� �����'�ުҤ���|Gg�VG[=�@��E�r���1�jΐ����-�D�{˴/8��+�P�o�
R�߷,?5��-C�%��2�KC}�&Q�bXC���H%�d�5!{��lCC*��u5g,�
��B��7��;i�Ll8
���W?�������o>tF�u	m�rr���;p9�ź�tK$lt�u�OE�J�c���4;��0�."z���d����C0k��W�)�\�=��W�Ș�,7Z�?�}kj�����lK�m�Yf�~�wz+��)���l��a�1�y��4���"�I��F)b�j��'�[�s׵W��`4��`� �Āq`��ϡ&������ݓBf�C���Ęh,��plY��5�[�7��7�U�Ep	���u�^'�]�S6���Ƈ�J�j �y��a����3�%&V)\ ^���O��~͑��L6N ˂�О6��*��@��ũaF�xϻ�?����Xm{׉��	C�w��9�;x��+�I�%7��|W��e���j+��j{xxI���Q{&�R�4��a��Ts&���2\u�a��y�FX�����o���z����7��Ψ)��U�)�4
��V���7��v��[�M�o��2�PQp���t�eO��SӦ��|;~̵B��_����a�'�g_���ΰ���2���	�bJ�t`�|����̑A�w+�ۃ8��l�U��4���)����Avu���?v�*�@�������f:* ��Lv���D�C��'I���tY�y§�6y��/�D��h	�*5�ƅCz`��`�(K^7��_�
���pep�#@-��.��O��轒.�M�VtJ6xǖ�}��*_4��[� �Ȫ�0��a����p0���sA�}���3����8�y% �.]W�9�*��G�/&�g�+e�&n,I��ۥ�#g?ԋi�l���w	���dM�Iу%��� �Y/�FJ��4ꍁK��������yt����>���8i�c�=�+�w*S�W1��P�1�O�@Br��g��SP+ihO��	e�B9^�1v^l����5�M �i16J#�Ʈ5�um��\L?\F	*��x"Ͱ�&$��@|��:�J ��u]��eB�ZQzŷ�Pb#~�+gj��`��@lL>A��uw��m���Wt�7�0�#%�_;�����]:��i�'���)�3)�e�
���4�r���^:����Wq�SjbG���M\=��e��X!C��+f��DY�+�޳���	�ZTN�;��AJ :3�G��EB*U"�����7��\
��e%�f�8y�������\��@��j��ĸm7嘒6��/]�$m
EK�8Hv�!��p�3�}���޶�
[16-�3�A���ZK_�
m�����G�Q�oH�X����7��IŠ��9M� �!�`���QS�]���G�����
��2�Y���k���1v]�KʽX f=O���x~2����N5��	bQj	�&c���$�������
��BV�[�\�N4�`�d��O6)�YS�n��/���n2��#��c��S�Bik���9TP���ub�n�,���W,�]P;��S�P��ͺ@�V��4T���7���̄�a���X�?�O$o푬V�>�
�q��ǒ7?]v|���L��e�df�M�p�����)����4�<�~���a�řK5�|�ʂX���:���('�7�q��-��ܧq��+"�u[sq`��5?1n�[�޻�Z#���9����s�&Y��rZ�����@��-=�'w�t��%�n��f��guB2ք'G�ʀ��MFD�>�)��c{o�nZ��i����_Z��6��s�8�	�~A!�z껸�Hy �va�wN�ò-�1��d���(�_л�汚N��svy��K�,d�8����Y�M�� �̏V�f��̦*�@�RJ��ƫ��j�??B���(]�B�d+:�֍Hdg�𔙦��w0uَ�5vJGN:�X
Ͽ@3;��_p�0���}��+�� ps^r�5&�g�܇�鍈�r�Zq�[!�����]T��J���|��d����.L�GF���,>APVꦖ [�x�Z�1� j���R�Gr1�n��E����*:��V�E�6��88Jqx��>�o	��ws�K����Z��;e8sL�Y��a��j�e������%e	w��RxM�V�l�����e��c�)���T���M\P/~����B����jVᆙ.|�6�	%�i�� ���W]t�K����d� �k�_�8Z�lIrF	��d��]`l��Fh���}
�k� �C�b��.��I��xA��j9�a����=��5��D�5��[}970�9�k�fW�X}8�)�+4�^WmZ��r�Vb�q��L��k	�@��01��$0���al�M�w�b��'e���'Z������fԱ������ڀZ{��K>N%4�xi8< 2OޤYә�Rx|�ô�x��Y���{YzFu�H��?��3L��Y�?hj��0��������?�rP}bґ�ޅ(��$�J2\��V�M���I''��T��<>	�hm˪Ș�=���-S7t����=&f�)ͼ�W��q��|�%��4C~iG��Eѓ��x����^�V�kW*J������('U�"�F��qE~��n������A3���aM��~��s,��D�K=��a��؁Spv�)69ކ�+5���{D�P,��Y?]/�p!f����ڸ���G����qsd�)LFy�s)Fv�H�M��m��0����J%L�-=�f�p�h䀺��W?pet&�I�DX�ϼ��f�s��Bb���gRS-�(	�K�+�1�xM<B��!i&9���V��������gBT�H�$�m����1i�|(��J�$�A�5V��]?�zu~^`<�/�K��eh%0���c�HoB�����Œ��Q���Jy��5�W�.}�	��ޙd?�˲?��)5��5f]�!k��� ��ME�T���>N0�\�1Z���CmԪ�� �[�;���xb-�GG���ݩl hc\��7�oC��q��_up�� �H7l@�um�'�B�ڭ��BLi�	~��Mm=�-k��)��ހ9��U6�L����u�u\�_vXL$;>h�(\��`U]�f �oP���K�yv]�l��Gv��*:��~���!AD�^��801� 笽�DE�>��f;�j�v�͞\D�\��f��LQ`M�\�m+Д"����k���� /�P��z<���?!��`��iX�k�@�Pn��eOTC��n�/$3Y��(xI�Hҭ�6Y�O,S���_V� ���K^
���z�R�}㴙:��{z}�PE�8/~ֆɪ����{4s�ĕm0�^�%8�`g�I�T����ڑ��X\<x�K���k YWQ�P�%��p��wM��d�rA����e:�,����RY5S�2�	��7������Պ* ~0n�dZ7�
P {�ea�mQ�Χ� �J��P4~��0y�:wSm%-�m�@;9��P�,����+O�2T�����U��'�Z��p54�8q9����6k'��WK!ۖ�S���!�٪�МS��v�oc�eB�w�d������
�DGJb�-������/1�h�rY�,�I⯺zuP�i��$�5�r
����D�ך�^s����t�5t������R�d!�E1� �wF�*:�;;E��{~���}�Hq�Y�� �-�@�A�*1ð�Ѯ�^�5��c3K��@��'������os�\$�4����Ǹ�1�(������lo�-5�,4u}T�����G��-V���I�X��G���&����anf#P���K;h̟g�}��;|����k�D�G�n��y����W��<� i��?��i2=��hg���Zs�����HG�as�o���)A"/�l���1��}���q��+�p>5���	z�pщ�fXZ"��3�Db8��G���N��ܯPX�4�Fa+w�ӈ�t^&|-����V��]���Uk]\���T�|�H˔Z���~�N�~�=Rpz�:�'�,��.����V�wJ��5���fԡ*,l���>�9��PI�ƥ	n����ԍ�
�6����zsx���b�1+cl�v�:����|a+�4��UN7�q��Q��WT`[������M�칹ޣ`'mE`! ��s����9����šYU�������%�|�n�5a�����7m���З@�qE�'7����]�p;pw�,�Zo�p�b��+|��qyb��<3lHЈ@�J�e��w���u�S\VK�e�V>����HC�2p�v]kv��_8􂲙�W��!�&}**ɸԘ�C��_��'Z�?��Ex�4!5��kRz�?n�`�Hu��˳��Q�#�v	�K,9m)r�Jx	A�2��a����ĕkw��Eމ�oA��J N�V�� ?��R�9����Q�[�������,Ý4��u���r����6�+�����?�r�g�\�Q}0�Rծ�F�%����fQ��+�,�0v�-�%SF_�V���
I8�)<"������YS2�� e%Ѭ8��U���S�_�FQP���=?���|E�byޓ`z��ux�a��-' =�/���NL��v�n�T���6]*<���,wא�+��<c"����~�^�J�@m.��H�r��×C0�Z���3_�?� ?�w̪��@Ch�KJ��Y1y�r\<��
���@����.�i%�cPM˫s�QĲ��
+\(���w�?�$�1��x��
Hm��I������	KN�\1y����7�����}��<��G��F^"���'��f8>Z̈́�^�G�1aa�D��-�Q�
k[u��lgԎ�)�S��*�*�b�;e��6���?�I�a.� ���2A��=_ރ��t.S��딝\�]�5�Z7
I�Isw�:��x��w|��~籃�=�L�(�6�omI��ey_(�K�?�>����������MP��7�]��@�����E��T��?Vն,?��+�����Bg�DԦ�j,F���u9���aKl��T���Vy�V�c���ۊCE[�2�bRaPI��Ȗ_c$8Z�uO��c�ޔ�&�TJ�.#�֩�Tom*X��������{�\a�|8��K1xjĠ�b��8�ĮU�đ�On���e��Z^P9<����;5��Ή�*,H���U�Q<z0���
� � ��8Q9�}-܌���QB) ��l��w�4 4�M��]��E��cծ��IoWtx ���+|��۱������0�r���X�%��e5 �waSC#�Ag��uf�|b���Ö�/�?���}H���ۆU��I�ѿ%�����|Y�P�+��|�hN׈��O�y�K|��/�sTo�gO�E@'�����Td(�(�b��p��Ⱥ�6�����+q�N�p�(<���۟���?)��_E�����Q�pû\�$e��&�E���D1=!���c
mN��@7�T���z�%���Q3�M����EVg�քUk�^DE���A�{�%�Ѐŋ:�؏�d�_��T-�Q��XՒ'��ʪQ���X4�%��e��i�i��W脭��_U}p9�Ue&[�u
����C�O����6��������n�S��S2L��*�^X���VжY�.��?��-��6�u �}�&��gꊥ�[�� Q!�2��������>��&�I�0hTLI륶�+�#��T�y_��qI��ھ1��X���z�bl@��NM���T���/����G8n���k�N��ุ�Oʡ�:q>����,�ޮ��إ�؝.ђ�w�m���H\Լp�g6�|�k���|\��uv��PT�.�p��R���lr׮����Zl���}�j�A���w�Ґ��jE���ao[���	��?I�E��5{/��[�N;(ո_�Q>T6>�%��T[#���|���܀�-S�O��]�Mٙ�	J��og1����23+Hr���`��������&�Ӛx�󧨲�MK1e�c�y�
�<7g��eO?V�#w���ƛ��L��lt��`q�߻�����0�Ro8��C3�ͪ���8���1��!	%�S3�i귄�z�L*Sb����ƭ��#b��𱒏�r�ܳr�7
3����y�0|����o�`�2���Eɖ���fj��Lr�K�&񒳯j�H3A����j8�mxb�I�MԻ�C�7GY��3
ð�Ŏ�� 
�|wj�S�A*�?����$�܂��Hk�(�P�f &�9��o���D���l���g��!U����Wۓ�,_B�#��jk�[#J&���3�T|��*���3�S��[ê6�����\�؃w�Pw�E]B��+!�-Zvv�9U�Hº�n��y���������)���0$��{˱C�Λu������8O�#s���B���A۸-�6t�읩���}�#�0��2�^GA�0�ipr1��o�Y#4=z@_D�,���FJe&|\��UZD����	=�$�ap~�dP��ci�U�[B%ۼQ��AjP'�g�:��;έ��]z/<��8� f��VG�D)Ԑ��TVC?)�{���5?on��;]�vY��V�{z8v��Y,�ksUP�lk��W�*�I��v(C֛�[����XV��ɣ�e�U������JqWX�Bf~��gtP�ͺ�_�VrMۛJ�~s�68���#ߧ�Cg\�Lh@}��@����0��/eQ}��9D��4�k�n����߆p��GP�L��K��`B}�c��C����AEĪ�i�L�+��P�����
$A��Ä$v��V1������`��{�{fح��4J�R�S����?����w���������}�oҼ�v(GG����!O��{��u!��ó���]q�NƔX��&T�'Y��}��1�$.�����_���_F�8��(T�A-�\�0���`����?͆���w�wɲ9
��������Ҙ��[ H^� )�2!���+������'��&���E1���k�c�7d|�1��m�tJ�g}�H��U�\T���,�A������CK��K������M�<�\�^+_ZAN�]�?ndr�8l��.��N�B�R7�#��QP<�5÷�~�Q��ɑ����ղ�`c�����u�(S%`T�
���������&v���%zX�֝K���j�	'��"^� ��w_}���_�ub�h�qc;�0��$�,���.�?��G�MbK��R�2y�maX����G\و��,�qZ��a� �-� 4��k6 `��̧
2=��8Hkm�9�� U͙l�F��]�}���˴#ȶ�]�bs����hkKɕ�4�BN�\B�2��}8)��&�u�|k�)n�s�5~Y
q��]�Í��;a5�Zۯ�ޯ����1���{�S�D���R,�/�� ���ɾ{�%h����u�D�֏Џ9��'P��� ~�\B��ά"e�'�%�Mnk���@<(����af���	���;���U3���k�S�P�$V�)B,�i\1��#UoC�c������+�UE��/���j��_GZ���g&�	��%f��tz��xf�ί)�)s��4�R�S/mr5c�R�N-Ã���s0���N�|/g
� �<�{��{:�4�7V�Uc��E(c����!�d� ��٢05����|��ǀ���o���P�o⋴p�I�F�N@�y��ȥ�=䫋 gW#1����Cϊ<��2.ֵM��1��\��kH������,�ɞ"?eyАj��Kg�)J���?(��B��s�m䭵*,S|�)zt��c�)B���P�c�W�����DI9��"�؀��7�PC�y!i4_���U�1R���#+�J'r3ءIA }�����"u@q�������q��9定���.��v^����I�������l��*��F��}�"�F�e*��R����$Yy���־>�ǹl�P��ʃKh�L藓r�e�D�� �����8MZ��KM��6��
���0�\�&Z3_�Ŭ��S���;Ex7O8P�c$o��䊀�9�6$:)�!�5P}^�l�� J�=��dR��S5�?�A�Rw�I��>'ҭo���U��Ne�Z�P��u��elk�˘v������jh��Y��Q�o'h�?���È�f�b1����^���Y��إ���)�nAK0�XK8	��-�W�p�?z�fg�8C!U��4��H���� H
��Aٙ� k���E$��R��/��<%�X4V��B��5�$��(��Ǔ
:���}VM����s�pH�������,��%u��`�/��f]�\=Ft�G�aL���֕I;����Ȥ	��"J2�؋�P�4��IcY��u�W����_��q��E��n�d���'R��j�pܴ9լi��Lb�S�=ںj�|����3U�����I�Dj�Kc���"��Lп�N��'�����*9�����L�@1��M9�K��H7��}ia�Vas����}{�1{,�Zė�r��BO��¡9��{J~TU��^�@����g��׎d�o~�ᡢ���d=�W����%UEo�}{?>3� � U��G֒��ȨZ[���
��=�+5�W˭r���Ń����o@ ����{��ֽ#���x��ʝ���zq3��hOށ)�E � �R ` ������U_��񣻶[d1~{�@]%Lf��q?�(���lյ��ez��1+Bx�/���sī��#�B��P�ZY�n�InG�÷T���(�͑����mݷ_9�&K��p���b�:�ź� �}�.I������kh����ƅȆz��["�c�A�(h��~) C�i�p�5OE�[�9���:M��e�|.w�{�ْ���Hv}s�8��KPe�K�AQ��曩�<N�h܌�����)y��u��+�e�3�s*�FcI�9��\	���,Ź�3ǜ�Q��%�>1��6������t��	p��8��r�@�|�oZ�F�0vk5�+e��q��6���M�?ްkӣn�gxa �����k�o����ā��gu#�q��J�r�����aV!f�Q��ր��ӡ ���=���C"�?F�S�;Ӹ	�e�w}r֓��16�O���Ӄ�@�(&aS�<��q�x�j^)V��;A��j_Il�V�Ei<=��#�%���8�36��&�]�R����[��F��H����5���J"��;�%j>�A��o�d���C�J��ɏ����sb���(��:W���e7y<ri���u�)��h���_��+��z�Ќ�?U���F����F�2OfZ�bb��<�cΖ�q����7��u��3���F.D���w��(@jf;�¼/iA�o�U�		��AZ,��g��z;;On*��Q�M)�s�\B=�odr�+�J`$^�x���Fx<�	�f�ƫ)0�R?߆�s�4ɗ�G;���?�Y:M�� `�����~QtH<��B�i�'{�l*.�d���u�5yE��
@� ?T���27����4�p���'���r2;�'����Q�~T�*�����a�Y.��-ǹ=%�0�!�V�
H/L��ޡ��)���b�����(�?�<T�)���A��,U�	Xd���VS;i�̞��4eG��\|���9��w����q��/�Y��.zԒ��"�B�Zz�oU�ɼg�1$� $�҄R�kwa�7�GY���Z����R���Q��Л��リ�A�2s�=p��c��26$*���ʌ".��،�쾫�Ф3���7���bH��^7��������\�E��'�OR�>n ��= �:p
�<ծ
�`An"�Af���?��D��Ĵ�VV� �ҽ�g%�,ҚUV��҄\t��9�Mڜ�@qr9=����܉f.���8l����r#S)�v�K���d�_=lAe����
��\<?D�<@��ZX��ŠV2�Fe�=M��2�Fgj=��8�`��g����O�!�KTTըr�+$�懙]}���-f-6 ��~��� #��5ϼB2K��W�Ui\`i�Y�o�9�����j�Q$m0��j�V&��A}bTT?�Zb��D�v�S$��D;�-�qM��(�~,� �;s�i7E3�1c�JT�sm࿚Wa��v�"�O���.ǋ���D�4�G�îl^�O�w�ʒ�z��0���]i%�~o�S�� ���~�ѥ��m.BP�/�UI�{_��U�{+[���j�9���V����x��Ŗ��&��Z
�7�:HB��#փ�E�y��=G�(����;�V|%C�=��Zz\��x�
t0PR��8����Mx�͑Ϩ#�E-�2�	������	�w��)!_���8���MJ4#�eB.W����:��3m�� ���ҭ�3@Yc��5�7Y�:r��Xs$9U���d3:Z鑦&�o3���\֑O,��!�`MyM�����L)A��S�5�����g:��<�
��_(Y�"�3�$0��O�)�]!"�`F\?\����MHL<�Ǻ?=Ý�_��D1���\�k��>�r��7�H�wo��c�?z����=��}�ryK�Fn��d#4���^���D�ml?��t<�>���-�U���Ւ��њ�+�����t�"x�O�Ɛ����#��M2z/M����$��L�t,��P��ҌUkM��g�Oϓ0pi��^$�tč�:|J2?!� �r�>�G �W�� d�&1?7P4���"����k4�Qɢ���0�=�VX����r֒�S5��^K~�%l"7�2���l/������nQmYgl����p^�bl`��[D%��Ȩi����	��Y8��V9 P��:�Qb7_1�t�y۲��}�m�OSbn���4�W�"��YIr��2�1�L+W��
8�r�)^H3�B�1V��-�f�"0����iOT����I�{�69��$�V����OP�Ȁ���ABp�N*��.-�X��+�G�Fܖ�w��- �"+3.E=MV�gL�$-j �B��;�&���ENK��G�>��N2�k=�͝=cC���8��c]v�\^x)U�S�^4����
b�����+�"x�����s��������>{\�A)U*ڤ����B���I��([�I9��h�'�v�������Zش?�d�Z�b[~�~��£6�R�IDG$% ۪L0������t�z<�^�2Aګmx u Ӏ� vp�X$Yg.MA�fF�7,�Ĭ|/2+;���)�T��'Badv���1��,^j�4�[�Ļ�n�!aa5p�O�_�+����?�6���B�a��9e��h �F*�-,��+�?���%j�P�����1z�V0B?�T�雠���6�~R���������Xǲ�&3�Uf�R�9�.1oZ�#�1"C��Z�"��I��4�:Zʥ	���5�����\���15�*�RR���.ޣt�:�ݝ8<���#�ƥ��A9��>��.��b�;sx��YlO�D�5e���-���$����M"�9������cHIi,���M	�9�ڌ��hc�V�t�����w���� �:�(w\�c�q�|~Ё$_��p�0k�Y��O��ғ򉤞��n"u�z;�.���6���y�W�I���8y�*ނt3��Fٮp��/ʆV⵻DM���v_����gU,�p �m�,��!��){��"�1A̪a�>�h���q�t�c�a+?}pm��i��)%%��#K�To?q�\�c��Ac%'��/Q��2`���/'�3b���L@=S�_���F���x%K0��^�SmS��O��t;��-k�� +����˶r����Cd7P�)H��9�e�t괖o�(�����:�$RgT��HM|G$��QCX��b�D�����?�C�Ɋ�)�#����A�]�U�t��w?�ձS��>,h���-v����z�;hD���r�?�R�Օ71��y�'���3x��Q��=�3�ӵ�i�Vm#��T�v��nI��JK��A� �Z 4?=��/a��}��zfs�ivd��tb?,���?g��mJ:�	Eң5G+j=�io���Mk2<�~E�>Fע�;L��3��d+V"R�Va�{�WmR޵�1��D�o�X_N�e�Z�}��@c^򼝮X��3��1�g��A���Xtc@��D��H�����P+����ڏ ��f/+I���1��?�p|�]��IZt`�i�\��H�D�x+7�g"'Me'l���Di�3�/�ҶM���J�\�X���Ј��o��q%'�e#�xG[�<����	���G<a�
uL��۠;�`ʞ�S�6͂@D�s�z>U
�����Ǫ@y�@�N%X��)/�.BB��H�v}�͔����;hN��>x�tjCQ+v8Ī����$�W�}>����p�!��X���kk�g_��X��K��$9��`V x|��T<w��сp5�f���Z�W��m£qŉt��$9��}t`���t�yL8h���ACO�C/����]]�lX��~`ܴ
/�Ɏ�N�,8���$��>�V�PM�d�W�$�h	r{���N%�F�xغ�Ͱ!��W1l-�^�ރ9�r�qnR�^�+� 	��[>�{���J�y�#!��,1�5Wng~�!H$|};@>��x��M��`"�!�WQ��2��jlRWKjGHie�c1��YH_��Oǘ��ΊK�h5j��Ze�
b[	[�ƌ�	�J�i蚏x�A����mv/ǖs�:@"Ņd�=g��wi�����y���AJh��ہ��d:]ؤ�b:�6i�6!�!���*����^�rf�6�+��iq�y�)�p��SQ���@��2�^����ܑv%Յұ!��'����o�z��$���^�D���_UU��n�oM@�z/����� �Y��.G�m��k珡�O��H��MG�[�&��3�It��l�X>�E����ہ���u>2|"�h'��
�i�-�K.D����0둡��hjTukl�7_y��`>�_X���Zz�j���ag; �W5����#G�U����aJ�0�h,;C.�D(_��68�H�$e}��m�B��C�KERdɤX�i_�F)|��8�Z��	��'6|u�	�۽u��|L��0��V�F���|�y�<C\	�ӕgg|f'!{��,�ȏ��֮du�P��DWa��$�V$���I�QW&����I�o��T�l���V��Z`���m����m�\��i[�/�
ފ�7��,ɝ�|�;���L�G�t
��m�s��*��6:O԰��i��qKP#|�9��0�c����2���7L+,��m:~I���x8��G�]pI7��c�'H��!X�{n��"� �/1�h� ���`��S2��)ׇW�:B4��d�@��PW�L��U/s�&&
x��=��TtQZ�����t"Mf�s�P�_�*{˱lJ���m�b��?}%���.��*��`�$ą��}ƺg�lJ�q��eh)t�]���܇�gqe��7�1s1�d�`�hhz�M �緑e��7����"��z��&j#d��d�S�#����i�/f���1��ê����#�=*��Y'�"C�j/7}��^���&�|����-"�J�d
pspsF�o����&|��k�P��nM�2�s/A"����8Ndj*��'��J��ܞ� ��j�R���X�$�0�R�2Dsny��TL�N-�%兩��\7)[Q@�/�N?����q����,k�{�cu���	@�
�w��A�� �����ruP%�C����~>b_Z�
��K�;ش�n�#|��%7OEU��"	�w3S/�_hl=�TsU�eF����,�E&W����P�l�) �ŴµD$��_�F�|�/�7t�#����Wc�l�[���EX��0�^���Zc虩ʬ�N3�?J`2�5��4��Ҹ{iCr�J[�8黛���G�<n�L�%a���F�9%	<��u����S�c����l6�;��;�$��O��B��uזd�Ek�V��:�s���Ԫ��)}���zy-0�9{�FI�E�A����ºkA^Q����ќ �nf�n��ĭW����g�GKɗn���:�v>]4���:=a��*�#.X�ݱវ"�jƴ�~�b��j�?�(􉦤����9�R$�� ���ވ�sR��?�������qg�+���8���L��oĚ��>hh���ֱ;��6Ay6�V��WNx�	~nH�ҩ�e���ܪe�a�ywRЄ�mq��ܸ>�����a1���dя�ݚ5b�^�|g,$�)���p����16�#`�����e£Fq�J�5;��������c��%�����s��TZx�/��9}�M;�Nw7�g���������k���7�x΀�fB�V��P����L]��a�Fh�b�r;,�&阂 a�� �R�!o6�s-:�k?8��|���|�gcB8�h2���)5 �~ma��i�O1Z�4*q�1"��i��S�#̻��DD��Xw�ү9�IxO\:�C���+8���`y�cݷ�:�}���Z,��*vzu����Ϣ��c-~6ވ	��tx��#[ܡ"�̵�<�Zw��x������T �3CT�R�(02�N�b���� ������^��۲ԿNd�lI�R��tR�Y+l�+�x��h>��{����?�'|��1�$f�1N�u��Ny��z-��gih�s>�HI��W\N���ts�ׁ�f ��Y�����>UI���z�Ϛ�G���
�~���s��~����cb/���m��+��B�T�2{�r�L�.��.�6��6�4o	��O�.�A��孹T��}�� �k��#������d�>��}¨��J�V�����6�pm��ZUAjچ`7�tr:�CB���K;�k���am@�/�";�1��K-�Ŷ�\�?��h��j�(�,����Y��|�2OS{ψ���y��l�|pq��oB�8ޚ�P(4�B����K�4Z�ՈM<�1���1e"�����5��6�,p>�ۿ�D~�i��zq�Wҙ�PTCW�������N-����O
����
4�e��dz	~Y�Ԗ�.G���X�5��ٍ�8|ú�T*W�eV7�d�L�R����Egg]].m �뱔*$����[�%c�ɀc��;}�Ӱ�������`aj)Ϟ$��,�w����*�t�\aR������JYi1�S#VΌ`�����$�׫��=J
o���6�m�|����_�Ѭ����r}��`��W޾�Wo�N�_& ��7Fȩ�F�u���`� {q����	5o�<��	��h�Cv%�_z�u�iP�P�E����+�{��}T��.���W`�G}-������-3;��ɝ=�WKku
	��"�S�1���$���F��M!��n'��+��?/6){%Ϟ9�(����Yv��"��n�>Ë�������D�ˇbH�`�;�vx��'��l��q��gG]i��P�� ��~<��0[��e.;����!��-$
��/`![/sZ�'� �����,������9��'@�{w(�i�����~�\ًH���Nӂ� 9� {�Ͷ�e��k�b�f�@���И*�a�,��sRb�&N��ŗ�Y,�$z�O������O�ǈz̒����|�eI�PCD.(' Z��Ϫ��z�T�>�:�G�s8Ѵ�[p_��8�,��64(��c�+�ҍ�5���p)��t�%��E�m?Q?�C	��w�����о������d S���
�4w ��8]/1ar�ێr�
v�8�W��gb�d�=��@�3Z������Vf>uI���ʔC�$�df~�YR(^Sh�ihR���o�ҍ�<� �S��N5X�0I��������-���귵�3v��yFV�*�_� gO�^�p�m�o����O� �l��FV�S���O%�Qi-��:g;�����i[�����;��2���T�)r�*���/ķ#k����7S�`������^,���ӭ�jn[TT>��"H|Fl�5�J�fgi���2���؛� o�ANO8rMtl������d#�c�&�x�T�JWf��?/I��(< �Յ�/�#�m�'�%�a@����DR��,��)ߝkd[Scg_a��64;}��i2�e:�ԁiթ�w�Gª=�s��}#ekv���'�07��ՑZ�n��x�L�����O�l���͢� ��*�O�����{�Bw����&�[�g�uzO���v��-�h�if���(g�+���a->|ZW�K:S�����_.��kb7�=���@T��^�΃Blf-�8��h;zȪ�D�Q���pl�DD+x�L��c�I�V���]o<d�y��w7�ͣVfzh?�� �:�J���.�+0����u㭔OB2&
v�YpDBҜ���e��@��Nx��nM2ER� ��͖��:��+��3p�wX$�Ho`f��t��s�xJ�c�Q�:9)�eP���C]c���-�_�"^\�+ �w�F�!c�z�ǿ��$���x��n��~Uyp��}��Q+.�@�+oդQ���0��S�A�6=�(��d���a��vכG"�É�%:��h��r�!"�v ��<.�x|TtF�s��Ps���l��t��pk�-n|�d��;��p1�֑�NNY����4z~\��J��E��y����z�B)8�g��n@��d%�b�W_/Nk���>��v��Nslb�;�Z�}�Ϳ��3����H*�e�8��8�I���F�g�w-֠�ɕS��хi�QL�Z?~���D|��$�iz��~���	��왝�y�_�:���Iz�ӟ�U�16�Zf�gIVkL�{�G�V�"={��Tn���%����c�XZ���H�_}�Ic���+V��回bƠY�?������V�ԓý�2�M���.%�2��Xh�R�}�1��M�urwh���#�T��l���	����̬^�5o��g\xL�j� �ɧU��Ά�*��Ϣ�]V(�?|��y=0O0�w���gJ��j�о���qS##��\�f?����Շc�`*%/. �=�զ�d��}� ���ӄ�J34���aE>�^��$+$[�R�޴��J�2}������xftnL3V��E�o2PX�Uڳ)5���:t�X(�� �0��Y�$���7f�nr����G)��SO:u��`��:�Qb�!Ii9[��9�ϗ���"0�c�a�D�Q�R鞹*(�������&��&|&�<�o-�	��/���'�$� ���>�Kt��]�_%z����������ye�P��\}L�$Ny���}A�k�#���	�oTO���-�\�)Cg��ñIw�7h�-	e!�Ab�T{��t-��u�u#��D�m�Ib�/f`_i*���[��	)n�P����vy(6�y:n\��xAI�/ŋD��e,ZL��nJg ��D/�<d������C=�GGY������(G*�t�Tu!��5���Ķ*���U��!,Ds�A�8�X�!mA��2Ļ�6X<�z��}Q)�+�@�Na���C/KN9rާ��
=u��|DK�TO�ܘ�X�B䵾�<�ݔ�c凪h#���ê�Mx�H��_,������k��|��2���Y"=&E�CD�O�O�|�l6t��%���g�pr�,��JW2p�df �Jt����#}#}k�!(���3j�Z�n������;�����)�)󻼭ƙ��Y
H�5c�c�kP,���Ŕ5�l�q��J�L� ��aMA;I�!�V�XvzЈ��d�&�I���,SՍ�L褤t�H݊.�7���l&��w݃h���L�ͣ%DW��\|��V1Q1��S8�p)���ϓK@n�!Љ��C�����P�bh��f���b�1��P�(Ȱ��`��ȕe���k[T���l�̾���l�(9<���jS�r�ϭ�0#LP�h�����U��tף)���R���� f�ò���+�y6��Wa������/�
7��U���a:\���-��u#��M�w715u�1����L��T�Q��<M���%��)�%>�(,��4=X����S��aO%�О.iɄr��� ���i���a�s��
��Q�,A�'�1���C�pRK�'�Ѐgxn�z�o(��K�m����4��y.i4f+��24Z���-�%�r���0���
,���.�eq<:#��$��p��Ӎ�.n�+�q��m�K����J���9rđu��j0��f��e\�YPyĨ��(B�N��
�`idl�"��hX������	�}h./ȇ�$��I���*�H.�#��߉\~B�G�a�h�.���jc��Y׼��$\�n�u�`T�8��W\gmլ9w0vA.TbCP�ˊt,4$�Nm��������?n�K3ʢ�p���d������%)����a�L5��X���zJ-'� Wt���/cc���hF�zk��R�s��ƀ����yޗ�)�r@����&����^�I��x��xr���?�'���Q�I�\wJ�2�^7(Y���'I[;��� ;P��< 9�x��ˌ�/=�������d�w�N��W.+ѡ�Q�M_�w^��;��`Zeop̑I����W*W�LX��
g7�b�>:�Q=ttS�Q�(۾� ��mH&���fk������MK����%��ϒ��ori5%�,b��N*��v���
|�8HXWd�ѵ��A<Nq���^7{��uޙ�`��ILJ��d��vU���GOKY�h<���u�Wv�P6a��h0�����`xZ.4��	�Z.�QNP@��i�fΓv��t6��Y�AF��Dd�#��ȁ���b���(V�����/�h��sI��5d2��&K'��3Z���<�KE���C��v���P-Z裳�"v�[��_��������2��2���F#�cן�f��o6��I�E�d�l���֐�щ�G�@o��r�螞4X8�������ﳣ���M��Z�٠�w&��sZ��1x��,FDg���I+P�� X���T+�)�e��a��>UI�0m��:N@�c@�X��,��"�� ձ�x�V�ϡ�ZN� �C�ktqH��tb�Oƹh��c���񚜩����`w�"|� %�Ǎ��2��M;[~;����G��ܗr6�AKke��Tx|tV´y
��\@�K
)�Yr9C҆�n3Di!�JS�;��*ѿ�t�iB>3c��`�ȸV�N-��E��Pmd(�=bYq*��m?��A�i6mbG���%�;O�@��QqZ����gc���SR���������#��3�&kg7í8^���>a�ء?R�y|7}�K��6^<�!�U�2����?/�7�C/�e���Q��(����M�����+q�^ց	L�܅���$��]�x�Q$�|<�5�"�z�e6��
n����Y�ek��+�L���i!��,t� j$<�ޙe�E��X��v%}��B��<r�g9$�2�v�7��l��
uV����9
4�"��¶�=V隔��B��ޥ�tμ�d[��S�s���B�/������^����e픞���'��3N�Y��C~d�O�;4���_Cޑ\�0�O�q������ޢ����\���c�(�n��j�H��A١'��&��+X�ѷ�0�S�� ���1��A�Ӟ�]�8��T� ��hEgd�zg.�I�����|��MW� ��<�XL]�:�
u+]�ݐ�<�-�L[VJ3TȎM��0�(:ľX#T��C�=3ۍ�XGQV���Q�?x�-y5T��
���,��I���Q4VO�7��ɊInq��Q��SE���e:'E�o��I� ]F���l;���"+����%�m٫�����2�}�v3�Mi,�޾	�BR�ĊǨ��7�1���6�p��F;�{������k��۞�����M,»y�ޚCĳ羍���w\;��=�!����D�Y��B^��13ߤqC���`�3�b�R�?5�f�*8�T>۔w�x��m���c��uғ���ɝ\	i6���
bYO1�m6�n�P����_�]{Q�~>�$W7qPS����A7����ia2���f�K�7T��܇�I� �/�C�#.��>�(hu>��i�yr{�B�3��d��S�%�V?��td��O�����o��dJp(j�����{�PH|���.d��'u�� �GG>�Ю��;����T�^��ptͽu���XY�����!|��~
��G(]̉��r�6�~&�{�ҳ��VJ�Ex�
V��ΖH������dL�p:n�y��%L�;��V���	��U��#��먝�4��Vƈ�㻿�o��m0�I��|8y��
f�ŚFc�N����Έ�\��]�� ���!v�走�5 �$6�չw#WD�J���J�m\J�.��& $#�=+��+�x��\{�}�
ᢣ��f��7쀬l�@��	hf_��`[>���3�����R7˥D���e�'w{z�*�@���_e4h
�ǘv�m�@"� ���`�=
b"��������?"��c�<\$U
��Ӏ��Z�/�+d�JE�u,K}߈&ƨ����Up��y�M[��S���uS<Z�9�-�^,�'���t�O� h5(M#�+&؅7�K�<DF 誨�,_�>�5���	�_� 9t_U�F`�$�;�+�@��`t|~�[���W�,�k�뱧�P�f=��r�mn�Ar,����r�S�_wJ@�>�S̀��}.�~,Q�)�I�yEV�����~]����4�ڹ�Z���+������{RE/�oX�.KQ�F1v���M����E�����i������Cx�Z��>]�(&��F=�ϖbϬM�*�\��8sdLؼE��,]��>=l_�'a-ߜ�X��}!��3�a�բs�s��Ǣ����b­���ћ������(D��K�	�	�F4��n}S��-�^�L����#�5gUc�X���.SD?J%:�t(A�7o��n�H�*;B���ԅ�j�CHF���t�g�'�ydl.����̯���Ejq�p2f�,Ps���K��^5����Ƿ��c�+�Z=�F͑抷8�|A��� ��%��O��~��|:Ƅp�·�nvυ��*���CC=9�|�;Ĭ�?��U_x|�&u���Jp z��I���dyY�pT��Y^�3���[8���t�S�a��j��IȋY�r`�����*<�7.�c�d|^tN�Լ����j��������"��Z��.�j��9K�GhN�rīP u�D��vD�ޟп��\�-7ؔ�!�$P埉��IQ��T�E4��4�P\X.�����dl�o������P�7��J�Q<	i���8:����q���.�{!���r|������H*;������밈s��jbh ����د/*���gk����PuxsH�%��J�oh�G�@"m�D3��W��4 ,Y/.��V�c�6 |z�Ϩ�@wMC>���u��A��,X��|�����7��lGmv�R��WOD�N.qf�i���7�^��f�C��{J�}e�7��e�[�<e���9�^j�i
v�̦mv9`Blb����ayt�v�q��ohmǚ�HpW�_���+����Fz*�����ڇ�wu��l۱j����g���;ʊ�1�ga�j�|v���|x�=�����" ��)�F�,���Zb�[dE謷�V�Tk����N�{J�鲅^���f5���GZ��J�j�T7��%z�9J# ��M��p�y����nv~{������څmd�F@l�j(1�#�Y�-��P :��2�j||+����~ܳYu��5���׌[�P�`�� o�N�#ԍ�؜;��9Flc�#W�J)Ǐ]N�?~BK��qZ}��v%���`ML����B��|�R��^�B�r�j	^�$A�)��/�	5����i�!���96&̩威o�ϖm�?��4_/ЌfM��}�h�.��F�c��"��M�}�{�#+�� TG�Ft�)ꪑ�d�O�-uz5*�!�Q�d��3�W��\cӂ� f�aA&S�܎��R6�+�y�{6CY~��~NƅUiH7�����O��<?��>m��S�Ɣ���:	��yI�|"�A}d�\�k�H���7�U���'F�`:���D򶇈�>���,�H�_ur�����ܾ��xK}��s��]�*(iv����'�h��HƗ籄@<�G
;j�"�W[�P"Δ؉��d����\9}\e��b�7{x�?gN���#B��8}2�F�e]��U��Ϧt�׌I���&�R�W���$�魣ߣ�����;.f�G&��RBo:bP���!>�ϫX׆5�r�S�G�9����m�FԆ�	X+�P��3R)�"�&S����iOH��a��7Q�.ɰDG-�G����%�ּ~k9�Y�}�<@�(�0�H�����6m��{۹�C���'��'f9����-�ϟ{�';<��)�#2��k����"�]M��~�ARR6��~��E��T�z�0�@�BV���M�v�h?���a��;V Q��-���hl��W�6J�����:������|-K�Ar]�[�L6���'.r��%��'F�� ������{ӃfJ�5"�����W��W}t��>����JV�-L�������Ĥ����*����'[
)h=7�ik��޷�!�_p��p�����vsd1qJY����ZS)��u�Ec��<_�Ŀ7]�Q[ ��rܐC]J�Z��p�+�sj��ܤ��R���۱�ZS: z��E`;�ygn��U~�o��_	�w40�-Y�0u�����
\ �ڲݿ	�dMR ������O,F�/҇��6ǳ�ҝ�c��d�������j���2����Cgu��S��l�w2���j��nW�ʌ G$�M|~�f4\����}u��AH��'ݗRצ�Fї��1�C�@���Бg�)��%0m^�>�V	Upk�Ţ~�3Z �P�u	��d��{���7ˤ�0��]��~�p���X�+\�(��
 ���P>է-��9�+x?2�p�ݠ���<�1�dU��'_j���j���-�D�էn�i��4�+��o�#@�Vq��8�ރ�HH��aY�lB1��g��i�vZ?���7��
崌�We��ޭ`����P�zH��,{�;��)8%��q
^���y#�U���Ċ�h �mK�L���|G���q�$�0]���C�0X�Et�:�0�*V�)f�h�{�r�����t�m�����.˿Ǎ�Q�v�e��A^�<mjG�_�7y���e�L3o�z��}�'�	���>��h�4�X�p�_ͼ�8�_JH������i� Pݼ�R�o�A��m��DJU��K�ܬ$��Rm&Sҿ���/Yŉ��#�Qe�����F�"�x�%3s�4�(�v���of`D��`�ͦb	��V" �c�Ʈ�7�q��҆H����AiU�" 40$��G��(�w�Wee���uL�(��o�Tϔ���Ϊx�)t����22a�� nj�tei��#�ҝ�h'H��+���W�5`;Kݦr���Ww���#�
x�0u����B-Z��b�wŌ��� ��Ѩ�l�{2���a��^۟&g�<Yɺ�K�0���j����9瘳�`��)9���X?������{^�!�<ã�^ǐ��<�����m*��5��;��ˍ�����ՀjW}v�D��` �X����*��#��gA$�5s֧@Cp��%��'s6�;/}�}�g��#�	<m�U��dZ:�+���A޺�!缭�ٚ%��z^ޫ��80d �������� �wV�6�T<؁B��<�N�7��M�`�p��S���q_A;G���X1����ߠȿ��PV֤L�O+��'�����'�d����:2����Bw$Z�Ե�X�COF�"S���P&lZ����W9��I�ڎ����>��<�Fq���5�
�%�O��X�h4�b{Cvw��;&{D��� ���A�� �z�%�#�{j�!�k��*Z�$<��&�Ţ���g1��������_W�:�m��)���&�
(����ī�5��ƌC�EзE/���D��q�7	�)�k���\!HN���cA���>`���I��w(U=G,%罎��x���������������`��N�A&�g#v�j�5s��<�� 䪗J��C��{�R�O���ܕ��7����a�}�b��XI�N�37u`�*������Ґ��o!c�|�D�[8�N����@_���п��Ō�F���ݐx�c$�mVN���c��&��S�/A�6#G L^$�)z��:yge#~���oҶr�l��֒-���O̺�b�q3����r殠�q��	�{O 4����n���WzN���*e��R���a��S׾�[��΀	�׎7�96X}��]Q��M/$p�й���h1[��H�ٕ�]�_��ĀX.�e;�O��BA����@�<���4-���?i��Vd/�_vE8��=xVufH��U�*����h�P��'�����)Xb�0���p�]X"N)�7C_�A�%C1jI�/�C"�}��';[�)����|� �k�J�M�	���a�$� �����4>}<	�k,�A� x��0�IG����];@����3��8�@&z͊�r>�y�V!���I[��gia/5k�-	K����vmM�a��T�[��E6{oF��>�]��_�{��˼���t�e��&�҉�	r�ba��Ejj�u�)!���i) �b��¾�W�����m�K&�c6س����hJ�(�����"�����*�7�G���f�F&�>&͐F2�:�DW����:��F����� _�Q��2)�ɕs�b�h�M�袃gVFQ5�=xja��������A�>b7+<�I�U4Ay��U�6���w�m����O"����>��ص�V�H�,�ҵ�NiW\)�ʥ�d��)�;Q�*ao��P=F}@�3����F����I�{�r���ls�	�bǳ�i�}:և�:�:
,b�C�l���HW�DA�Zځ��ӛ�̴]��HS�fL���|%����L�����b��W��V�[�@͓w���a^j�Rcq����}�ۤ?�B����y�{��vZ���j�ڰȫ���~�V����%�i�Š9�nI�.��5�f9�-+c���{ܪ��
t�P@�Ͳ�5�i'��iM� �C�Q�����-�p_�ƃ
Zh<pͪ����Z�j������}�O����>���.�3��@�iY��K�[�����>��s��=1B��u,i 2F�n��m�cS዇�E70��/(+`sӗ�2�g�^�"���D�o(:������+�b\$u�~w��&�r���x�����~�(���{qP�O��s��`f��7�c��]r��Jt>�������u���p[_�K��	jC��c�f&��иS���ҵ����\p�ܢ�/�V��S��Q�R�ɿj�� �>���|Af�X[��ٶ���0�N��D	{F�]5��-���:�[0�	(���k��:\ۂ�{>b�BX��?�?�u��Or� 7x��h�=������Q*���6�L�"OO�~k���>�� vޘ
a��t��Ռ��ƚ�<��B���?{��?��<�1�Vϙڐ7ly�������N�� *:`�V1��*Wj �F0�1u1����۝��0��u/t��o��Ȃ�&vboL�vH
�� �K���'}ܿ��^�2�7+�6�K7Ռo���$#U����WbZ��j@>�����"��{kI���"aOqW�䬔�$���wT�l!Q��Z��0 �O��G=]�>'�����Е���GŞ;��J�UR�P]����v3+]�/a�)��-p�쩽�3 �;�y-_�r�o+hr���S��δu�� �w�/߶��)MoJ��q��x�������O��|�B?ٕ[Јm,N1�&�������b���'���q�5�������%@����oX�X=m�bs���`aV���[{gn��N.��"-9�+�[X�]��ۊ��v�HTn�4���ʙ���js�E��|D^;����bĀN��s��/���y/7�-N��?���<�.��}�듷g��N�J�X�{!�����[�����Fx�&c7 K`�/0��ʼ�x4��z6�W�9���b����Z����3�����c�V��� �^���_'|��%��_h�
9B��<xT�k۳2^���+g�qng"ץS��>�?{�`��Y�������2������X�N� �7Q������FV��@�n�F���9���P��u���� Q�- ,{K%7⪉Op�����$9Ez��QZi�F)��L�ݬ.��Z7k��yV�a�q��9E�KY���X ��tuab�O!��b�HjB��c�E!�2HE�}���˱8��P5�f��|��SSo����.~�`�/��[[��/9������菥���UGi}4lMD~��
�x�+p*3��vĳS�pf�|���������c��-č�ݵxِ�kg:w/G��N
�T���K�TM<��qjM��>�^C�k��y��Tb���Z���8�/QZ�[Kar�Ȇ�e=4��u���mǟ-[��G��o|�l����YR�g�f�C�GX=ߔr�N���l����쑩xq��ǒ*E�����KaVN=����6z\?ퟰ�"hc������E�8���)ZEͿ�����0���]���0�cl?O�>��(���{��
e��9��+S���X~A �[��.�^P ~S3a��@6�����r�3�+A�[qN#l��.��_g��7}(c��:U�i`X��1�8;{Hx�؏:��xr�l�h	��;U���>�i����A!1v5����R��4딂S�Fu�g���EQ�4�>ݰ<O�� �c��
��9.�>���4�Ɏ~%�|ĵ!T�$�6޸��l����1�Mv���Px�1�y�EZL�a�����H�zȰ �6�`��9~m�'���z���u*���0o?��-5JR�m�l
 ��^DUn;?�`�����>_Ed2C��ʾ�0)H�p��'��^z�L�%�0��ؾ,K����@�N�1�3�edc��DDZ�K�8��>e�8�f��K�w�&�y��F��"v�T���՟��ƍ�-�_k0�T��&~H�����я�ά��9�4r.��w�6%bR��l�c�s7��?�d����
�~�[-P�@"��֤As�E�;�QO�_\���e���u���`:z����:HO �\�k�/E<{�5#�B�Zg�d[Ի��3��gZ�k�Q�KI��Ȋ^�9oڶ6J[�-r���2">��q��3��;Z��HU����vw�����n��=��^��A�7����ǩm�f���"> jħ�sN9S(K_�&L�n������8��K�$(ҁ2�iی$��Bg�|�)���u�r�0xu]A�
3ߌ�L��[�u#�F��ݑs+�K+�N��u��b�$u��X]�`ᫎi�6_Z!�fc�N�� r�]ƙ�V�'��F$G_� �,CP&ܪ���6���	ʌ��6n��v�>�LG����>^��}S�!��&�1��d�Hic�Z���k�Q�	�8z��g���lY�S�Zo�S�6�h��������V��)h��JF0(mOġ�22���Ny�J�:��Zc+R�r�!�c95�0?J�Ofo�$�qV�R)')�O���tk�w�`�Z�<R��y�E
��u���YCy��t�e�h�����fT����F�L�t� ��dd��+�u$�I0�}�q��e�W2�(��h���'��_��57+�Τ�`�ga�'WU+-�� �Ǖi:\��<)'���}��ZL���	�G�T$���OZ�4�o�p�d�y}�A����Z���Յ������X�O~�f�I!i��vVuX��Q���L1)t{_�NG���+6\l2�26��́��9𪜎�^�����U�c�'�86B�.�O��`��Q�$w��1��hW�#��>�����Ɲ^�Č��q�ⴆ	B���M�q����mVo�&�Zk�I��Lz´�D5%^��`ӷ����d����*�``I �-� IS��/�ʦ=���no�5D�y5+���qD�(;���wH��Q�seF�j�p(�`d:"�v�NY���!�	sM����=X��r~:!�8�}�����s%�mF�?�X�:-�{N��t���q���*B�F��k{6��O&i���odS��^\�޽�X;��T�kT�[9��U�Cqm���
�zS��c.ٸ�}p^�}�K4��+*��cW�>��3�~��/e��ߞ�湚�<q���.�{+����H�oէ�[9
H�$�*�7�N��C�1g������%)d_�����	L��H�W���6����BY�9�ᤂ��ϩ��_����IܧM� k��4Գ���+��k>�k-.�Ux;v`�K�≴���ŏ9򇞪��*'�$=}L�.YZ���,7��w8�kB��� Jh/��)���p��j�|�oeP�2�D�D0壢�Z�0���8��9D:���j�w�iZ�c�\v��LTL�s�/X�DV�6^�M�O�����ȼ�>�^���9���!i���N�ibܼ;G�V���PS�!�ɡIR�G�eX��&�q��u-:q�U��	GMMN����;��k0�Uej�Fٹ�ހ+���[ȭ��泃s���1ن�@�7�&V����wDH�"�Nn�R	�6_�F�:�ٮ!�7������q7h$-��n�K�l��ø�[��K��D��Aq�X��=`G}�����V8�2�I��נFDp�$��P�8L�g/V	������^�{�Ӷ�^=�z�N���3[�b�,�i�0�!95����r�S�300���x2�61�gm�j�9c�|q��ݼc	�@�K�K��Ӫ�d���@F�Y�� ڐ
�L��������}��L��b�/�f)KF��Q�g)B�Mp��)�*b��E.fD�?Ab��G�z~���(�g�yB��5һ�kJi�9�X�ܬpx�HTh��m��(����k��F���t�g郐��XS>+�rCH�w�	,���L�6i��%�b����}�-N�d��#��8������r�6�cz��b��,I��:<Ϗ	�a�W!Ov$��Q�O2����Xl9͑ex�v�fO��-c7��)�����Q9�HSγ�49�J�n�ڂH߯���3 �l
�؇i��¾xd�����s�/}�d�K�<�����f��;ܪ&�e�M9e]q�c��V��)�e�d�o�N�<ܷ>yf�Yv�:��\)>�F(��
��j7W>�Of/�B��d`$Q�û;C�)ci��P�"�{R�C�9|��eȀф�Kg!F_�tӚl&�j�9dƖP�%��7bT����/�c�@T�%�EU�`ծ�b���t��b�����NzL�¿�j�m�/ĐU��E�I�#wcw�~�Zmr��f[���f`ߊ��;:V�j�w����4�ʑ"--	��?����VF���a��O�#9����OG.�����,l��C�`�����m
�f����������4��m[,s���For�+�7�L�]�9?��7dI���-�M!������&F�'͛wE̵
���J��k�(�u��"�#a@�t��U�/F�ʪ�����1r�/j�)�C�����R2�ٜ?&���IoO@ׅ}��U�t1����� ���x�����空��8Bb�L�>��\.%��0.��g�֤��L�;���Q��ܳk*�����Ik"c�������u*�0;AE��sH��ٕ��~��p���� ϞՏ�;���<�,��"{�����m�%bf���[+0ߌ։����
���W�︣g�}����}�B��%z��Y1mV���9�?|��uN�x�	f�ߦ(g����Өl
�1s��5����5�*�~6��܂�w�h^Մ0�������Lf�;��d�B	��s
+�p�8II86�GU6��K,岒OC�g�!b��4��R�q4,�1�cIYB�&C��"�a}g%d6�҄,!����V����\���"���u�Ɣ�wǴ|ʖ���<2f��<a����e�*��hf C����gr[��*g�@��&m�q}`N<Q�f�.��&d[.��ѺpB{��mx�Q��>[��wqr����i4,9_1]��H��H0���p<������-_{Q��[��u��.򖧆 �k��uT��#`�oE�-�囬�Y�V]���HP%�?}�����5���^��?g�Fc�����q����(5���Z�ȭ�`�M�&Pm���9zu�]�T��g�d��|��GNTN�3e��%��#a����m��L�_��-a�d(���.����%ցܨ0�nM��Ť;)� �o�b�!s�� Y�h�:�U����!&<�.�	 �t��XgÞi�B�a_����%�Q7��"!`#6�N3�˿��O:_m��j�$ۓ�L9k�����ˣB>"�kB`�Z�ؒ&4����qv"���vL�.���MwȖA�Dw���[^�AG~*�_{�i�}�~\�LGn�Y��o�Y��.u3����-ᘬ�7�YR���^��i��
��<�k�������b/@�AG���wr�( ~MyP�;�]�;�������8�\��2�l���)^��
j>�0=���,Z�5������эm�إ�%�GV��oa�n6JҚ�jϜ�a,o���?�
��:�J��L��
B�1�7�oQ��#ryG��K�t�ta��S���X��n��s�ڍث�>���Vg������g��/��&�%"A�[�B�n��y��j"@r��Ŋ�D��!slw����$�����x��.]��^�pJ�L��4���ǵЈ���.����=(��t��D$��(��83���=�
��E|R|KәMס���1p�$�Ѹ���_����<��śt�Q����&	�<����SD�ƨ�� X�=cv�~��P:������� ��2c��~dtXI�`9�b0���T�kɼT=�`z�/�3 gdV�XH���|�`u, �Q�E
�:����!�p��lr+a�p"��؉K��X�r�b=�h��^v��&mJ��l���QBP<{dA��$�SO[p
�FWW���H����DmF^%�5i�t7cW���j�����{M���$��;"Vယ�$K��~�I��7j��S�E4��Q?��ڱ�:����x���"��;�k��j�`��K�}�M�L��R��v��w:��O?w��z �,�Bs�w��pO�=kS`&iu��(�n��ֺ���]I��x��-�X�:
�)2�����@a�6������������,Y[*�j��;ym ��}?FnT�p�cЁ�uy8z�?~1�u�XB�.d�Y$q�����p��M�i|e��\M���&�
lSٷ3{��:oBc���|_lfY���Ix�Ya}��������_��ot~�z�B_��8�P�Ƃ��n�٧�a��JQ���2>2@����lT߅���(��'͸�כ�2���}�q`Sb��zM+�F�ߺŘ�2a��f�^�/�v Ul�$��m�8,�^�}MMB���?����|��Zs��J�Ê�a2�3v���B?�q�$�����3����^�=+ I�$��^q������zϸ��	+�?��
^)^9b�5$��h�j���0�����`~���_$C��"�ؑ&J'gڛv7��.�_�!�I����[������I��e]t��mC��uЎ�{R���b��-�fU[�A�����FN�X�B#M>2�:�5�_
H %!��s(��@�l��"�A#=X;��Ί����x?���	$c]����L�	�>�ś���;zÒs���?�b����!�_e��r}�	�;��iJ(kx� z��)�"�Z�޿�ڃ-�sD�wN�(��z�-T��Fa��s���t).�Xǃ�"�~QK�ʒ�Eo��	*��D��J/)⅃��{�4�z�����HIaP1�=C�I0��AH��Ξ?F�2*���7�UM���*�q��ȞÀ{n���s�o�k��r���K�ч_C���O�lS�~�x�z`���g�����̸!x����}~�!� �@��̎J�M��lb�|�e"�����eX��l����A�����j$Tv&�͂���*��k��S�i��p�O{@����a��]�����c���� {C���3�DG��J}O�>�]O_�����1���2"�Ls�m��3�A�T���0��7�r��O����%eH�"L�z`m�F2�d;Fj!��ؕ����#���b�՘��M.X[� �D�z�.8�k�gLXe����e�̷����5=��� �2t=Y���VG)�}�W����R􋘆1�'b���fˈt�؛A�����~��I�����ץ���˖U�0�p?.��tn7{A˸���|��\:�rq;�/���Y�<o��`X�'D5̪s�'a%�t��<����y�f�0�uH�@���>Em�_W���` nz"f��^tSA��&������-��T���	}��n�$���mY���Y�U{���%�jQGf: �'��E6�.�
S4�exo3�[i8�L��̍Æ�e(Iԡ�w/��;F��z�N�صf]ϳ��TvB���zVl�Ʌ?����ߜ<�e!E�|gd�Dh�� ��:/ �p��Xy���%�~���1�Ͻ?,�$w��EwJ�=NqU=�
'J�;y���O	�hy�/A�����/c[���u&!ե#D���:�4��V�B�`�p�5"\YI�S�#���K����R�fŤQ`l��Q��xt��~����%䡉d��s�9��4������u�j	�l���l�c}<�s}Re�v�����Ѯ��3�$(zlUv�W�w˗M�:�fH�'F����@��'�^Ox�@����	؎�s���ZD���5}��&��2�;̗)�|>�R~y	ߤH�_=D�ђ��fX�ں��8f�@ ����������xK� 	�:R��q_[?P�V�]4.�7�j��h�wp�3�Q�8�Ϩ���8>vꖟ��#��������,Bv�b��d	ǲ�K�'h>kqy~�i��o;�o�M�Y�¨��,>����dn~��8�K��DMj�v�}��ҕ �Ҕ�%�ժz+�Y�N�%�8�3���G�v�Ӵ�sX#gWX(�������w� ���/��O�c��F笱�c�Z�/�H]4L
�nۓ����ĳY�(Q����I��r��9"�Xu^탏�`!���[�UPC�h񍢋��Paa��cN���&gf��c[���$�>�VS��}��UX�?Dc)���sz�� ��?s+���5T�����F
�1��]���`�E]_)e���@�Z��7^_���=���kE�y����Q9*|��q����PxZDi��6	�����	4��)\a~[;��@f;���_!-��V���y[��J�ɦ��P>kͧȂ���1�9+2M�6Mq��7����A( ����MB�|Ʈa����H�n��}��;3�B��/�}BX�S�)Ӫ�'&��nvE�k��- �������mPY�t	��)m������+��Y��WRM��^O���@����M����gK6���]sqߘ���	�0��	N��݀ʽ�d�T���c��`���-x@�h3����'tm�����n�E�h�L�υ�|��?�hK�b����n�6���o�6C|$���Э�]3�E�%D��$�L��8���j�	N#<@�3���
M$m���Nz�v�����>nI#}����K�Ň)x� ��Mg09���-�?x�Gr=��2��=WXiZ��D���M�p���}������4�0���V��U�a� �fʌ��m�ZnE͖`y��f�yaP����=�F(`4&5ux��|M�w3�'�o����X�Ae�4�	�H+���R4� �0�tij�h�5"�]��3�w�`\͏�m�i�1ȿ�U)s:	���)����!�'�]��p��8!�a�dx5��Q<��-��r��*��傩���|�&�}�fV��N+a�U}!�y���u�H/�Ų��>$Vh�B'�T��
jև9�Q���,vRSs�a?�8���`��򳰘Uy��L@ ����>=�����;�P�z�Pg�t��1Bg�����%�	$k.q\�o���k�͹�,�X�MI?����*��zy�E7���J�x��vi��`v���<���Pu��z����ġ����r?3���Q��8����-,���^І�|8�Vw�����3��|��M��Ɇ�^�le��0�![���z�����~�i%Ģ�J���2*���v2��EPW��%񆴨�H'�5N@x��$������p��T�yc=�a.���>A�"���E�|r���0�Ѡ�6�f!m���)n��e"�_E��4HN�Tw��}� j�F
F��oK+���C wR>��/�_4��dpO�5ټ���7�:Vb4�[�-Z����W��\"���7=�a�4v^��ߠɨw�F���*�@]�*��!����܁-$�.`��`��?�s�<���9��F��{�9�Y�k��(����S�c�po�z�=]�#�Mk�k�J�)�{Z����V �ߌ�+���C�GJ��@�RR�9�&�Y.��^���4��J:�c
���Av��_h+��B�nǴA�n��T׊H�E��xэ8��R�YN)��f�ߙ��
��S��\S0���2�`�B":�8�� A�De "pBlm Q�鎭�q��:�=%�#T��9*��Bg����޸�,�g3HSZ�
b˴J�e$M���������[RƼ$��:#��4���2I̘�U�#�Z���>�)c����CC�F�x��˨�x����*��}ppH\�H�=J	G����AQ���V,U!���OՎ�nK��r�����!Gq�(:���%#]"��\��T�tO��/)��p��
*�)����iYIx�����F���r�ҥ�	L�&�i�~l<bͼ��������ׯ6]Ȣ��o=�Sk�|3�o�������'yml��0ډ7~�6*�9->�˱��ڛx<��o����W�JM���jU��X�Mj��bO�m�:F|�P��â��q���\@���]�X�-�ɳ�Bs�F�s��66/�Pz z$W�6v>$M��r�'��	M��0lUF�Թ���S1��eW� ��?!<�7V�q_b�S�| @|�|˞qo��� �����
�D� � 5�����x���7*��h0�~2$�i�dyB*H�'���Uj��D5"G���A�h�;�I�a-XR�����@ea�=�]e^!*�Ȃk��|<����O��uG(M��8c���´�.vג��QsP�����r������ms~�ߦ�G��V��I<����\�d������z�����W^�vi�T���vu��LU���ɲW�M��=�f�9��m�bl}�2Z޽����+	lvPˈ5���9cU��L���gɗ_�饏����ЉS��7�lV��Q:�U�� \�S;�ޝbm��t0}��̿�v3�$6�l�}@뷾%l��C�C����m�#R:��tY��3��P�yo_J��b�	mK-�� ��u�Z�O�P��@����{�T�mⱘ�:�q��0u;/bR��M�h�m˕�0G�E�Z�����u�5	a��S��Y�Q �Jͅ�|�mD��4�)�g0x�]���-��(��0�N-l���9eq�����<��ө^u��!;2��8�-�ܤ&Yw	#������۬
��;�B�@���������@#�N�&�J�h|7d`�j�&�$m��:�����B&�xR0�/��$��H�m�����& �xy�D%����#��4@�>���^N|�drv���[4���q@E�l�u�I��%��D�o�r�s+t=e҉��g..��uM��#�F,�޺8/p�I�p���� "=*K��x^5]�@XKN|�T�J�@���U-@6�(̿�o�=��.h�sÝz=�ȗ�Fx �f�<�k�;(�|fD;(�h�g������R�J\�J��A�?]��Vb��E����������������(B���$�$8|�'M�+�s��qwS�����v��>'���W?�vy-�S�2 8�;2� ����d�:����v�4��X���W}k��2����.Nа4
G�[۹o�3��v9�̕�|�5�������#�G�LґZd�g�=���W��AY;2���|"K���I�nc;'R�#�'��W��?�ũh����t6]��vڣX��H�P���Bg��\�\ȂK�!����
 �ə䢯����aS�H���!�����*��ȩ�^���ƒ��D��k{1M`}�#P	2�͕,�o�H�{�	���rb�Ƴ��6¿c���|<n�Qϔ���Ex��t����0ؽS( �fR��w���x�j�M�c�>0znt@@*MG����o��9��ĜC7�$�1\	�$19��؆ʞt�?�A	�(����§�'�Q�L����0+k5	/�,��N`=��������|�@��������	s86[�G���{kG�G��N��薐���Z|/���ؾ/ܠxX��ט�M�> 8�v5�\�W!1y��3`X������74YE�]�u8��3���C!�5=�љvc��
'��6<Z����w���?���v?����>���3�m�o,��`ur�a���%Q/��tO���V��e_��J]�h{_�#/�L���P�"ۺQ�h�_�B��`�y�~�#���/����x�5�kX�����w��gq�%��6�H3,����X��Rߠo�G<�>��t���W�?����R޻�B���c�� 1��?�R�vK�s�
�9(�N�٫EF	��׮ ���;V��Yq��z��D��� �2W�nMb��n�sj�q߬�F��/cR��C)y��V���ZHX�L�����S����!W��v�\��!��G�X��_�����\����"j�8���J�s�ټ��N�b]�A'%n��:����
��6}���/�ƦD�f����Ċ
�4�'d�t8-��TeY��?�*]������$�^�U2�V����6�>����l�L,$��@=H���w���&07a���,ڿ�ǾY'a� �f��ۯ��6��~AX�heS����4�$���"=��l%|�M�Bm0�W-!a͎U�:��b�"�',Z6��
YF
�^C�H�?��pBIo�>�u4x�q��:�E葭Gpf�F:eDFF��C�*{¥���í�����?w��f�΍��;�Af�8�4���(o�yCK��SU^��Da޵��(oH~����Ŧ|�l[��0^a����-.ъ�n�Ngk���'T��Pɫߨٟr�+��G44"��:� �+���恔�:x)F�н�`��>��(�*?��2�c{5�Ȇk�iksחX��w�\%��x#?6K�: ���I��P�^7{��%0k�Q&�����O��L�-	7�1�x:�����Ћ>�n��_2��7ȣL�
ؿ�$ 0X�{˱%zJu���;�,U(d�{Ml�v���D'ܢ���p����<!ZNh ����Ɔ�;�㭛jwz��`M�[Ռ�hѸnw��$ 'Q�Ϊ�g��v/��@߆+���ś.��a���=8e<�Xv�8{BnA.V�x��l?�t��\bE�y��:{�X�y[jW��ʎk��5��mw�����'��훭(n��H�!lG�|W�y�}�aJi�h����b���
w}���Al����ĭ)�k�Y��/����w��vY��9�B�U�$���b+����l��ӡ����2�<�3��Ӵ�u�%D\�k_9�Ħ*H��D*�~���E�G7�C�?=��)Ë����x���-��1P����ǍXp���?Mb��i1�ev�Oi�.�}�?w2��(���\���>w��+q��B�օ�#-Y�e�����d���^`�sZ���fr帗����j���f�4���Tv��`��D�\_W)�C���L�6Q�7b��M�a<u�~#��^���[[:�/U@��s���\^w7	�E�k������@[�����S���ع�);/�j�Ms<�O�w<�C�I>(@.UQR}t(P]v8})�㹎��8�c&RS��^Ӥ[mtj�J�C���e��*��z7�%m��"_�3��ۃ�	�ڦ�^��&���XԼQ�x�C�Aܐ\��C��S	�E�"#�`����BH�w�*m^%��ss]d��JFBY'��"X��	/�J,+����wok�g�*�s��]0 8l�B��S���=7�ڠ�{�y��#.ޜ[d?P������SB�&�?�H�T�ͦ`G���x�ln{O�J pMUJ�|�uq@y�ףU�R�5�!;����p�Zێ+��<;]6 L��Q�����:�e�ޯ�eAKs�l12�~Q.T�ew*j�nm�>�s�|[04�I����@\�e���0��ԚU���9�,�&ﯠp+���~u9J	�U(�
k�E�ԕ�7*!T����؃:ZL�c+�F�`���4�8�3Cj �|���v��^M�:���~�<RDB�u���./r��|��Q7x���Ty%5��y��ɱ�`&���r��uI?>൩*���� fE��6ĉ��;�.a�j�T��j5rTzá.\��PԻۦ̴��8�:�>a�8{��$r*�C�|O���_%���˿�nw��s%��A>S�*nma��6�R~��RX�2��I{�R`G�	�p���O�<��_g�!�2��iGD̏J`�]_
���O���T�1�� �3e05._������	� �+���D�_0�eg]��"7U1����i�;A�����+8q�(���S��'8���b���'��C�(����^�w	'#�C�`�n
<�X0$l�Du\�,F����oV��XAP��"�����+J+��{�l4!vQT�y��D�gE�N�l�ʕ���{lXo �����̏9U��;�T��i�%.�L��rP�aE�N�)�Bƥ�����*Z-���K�ǔS�@�3��dg�/���u�	ˤ酇E�,H#�R�"�dh��\ y��L���X{e���Y�w�E^���9�Y����ER�gX\Wg<�Q;�ӏ;H_<� �%����u��0Ul��/���s���n{�ǂeٚE+�9@44�ty��z��z�I�{���٨�����7S�`:o�:�a�%��9��i�H~(��Մ�U��;L��#���J��̞k����
��M�2z�?C&��#�����?�����"Iu��������cze�d�I4s�w5��d�Jm�g����"k�8�=�>?$��i*�N�#�x~*�Q"&
F�^X��Og�D[��o���w�o�9�h�J8Y�Z���]A7�W�mi�&K���h*j���2��� �XW�.a�7;&�8���lu�]U��E���y�]}����� ��y#�&$�(f�\&��	C���6�#����{pr�L<7���G�%Ĉ�[�
�g-֊a�'��U���"�����b�(��%q՜��SfIZ��%\!wq_��P�����k0�������V(p��j��:R�M}�k�]�y&p�T����l�IM�5s�ɇ�<G�Җ�2����o����Jm�Ɩ�Q�:R�:κ=��FfցP^*R���+t��@1/��1����v�~�~
��b��?�:'Q1�
}���Z�B�S�WD4L�Oa���G���Y,��Uf�S�ep�η$?�L��p���yʪ�or���v����~`�+��n���7�Hd|��l �7��f�
�ꯀ��c���H��7Vx*`"o:��)3�:�r֪h�}�����ǣ��>����hLb�	-*��:���~j�R0�x�r�FPm��������Er4d(M��1��\n0�g�x4��z�Y	Xg��8��I�!���O�Ty����:*WJ���U�_㤷�I
�JZbnN�q�I)�{��G����	v�#z��vpY:���ƀ�1%Us�������n�*�A_F\C��Mpⴈ߹��"06�+&�-"P>2Y��8���oܩp`NαA6�/F�+%��s�G�Czo��6�k��qk扅��+�3P���� ecG�bZ<�F��\	���BROy��'/D��Q�x۸��(LL�qM(�ţ7���M�������B�����Po4���_�л�r�zD��0�.P�N��-�*�*"�u�8�����
q{¨ʤd����D�1(&0��G��p.�m��9�i�2V�oq����8�N��9|%��f:�LF�4��k�o ��� ��-:f�#��"�A��{@m��P٠�����	gE�)��[�*+[�dD�$x�6un  oIT6�\�w�@��Sn�{@asQ@Wܵ1T4i8[�fk���JJ�mp�iJ�9�~m�
=�v����
�����D5�n_����{�Mx�J��K��U��Y3exQ��/O�����i�8.�,��,�f�@��%���cD����I���ۣ�H�
ra�I���r����^܅A2?�=T �4 S���T��2�1�ՄRe�N�r���OH��͒&��\���X�\t�|��lx֕SwJ�X���b�Shuhi���y��	u�/e����2�;��H[�,V'+�;�1B ����{̳�{�=��
�ش_-��64�Bs7�7v^,����z�qժi$`�ߴ�q��Z��R����Ռ�p�� ?��7��(U�x����/�F��s@c6ޟU>p�=џv��I�4~Yl��n�>ص�f��MC���]� q����LLfX���f�%%��9�uu�&y��鏌�xUa���˫vЎ�2Ft����'^���C�B	�\/� �}��6 ��&i�3�m��,C���K����Ē�9���<�� y*�G�N�P����X[��q �J"����z~֥�BʱG̍Th�(��h/]�ĒPg�o���=��@ h���v�	b�y�B����d_�k�f��!��o�����Ҹ��������P�3-]5(�H:%�o��T��yL�2����Y�W�(�.]f�i2,��(Fk�x�.�g���o�{D�\�1��"��L�UI��8cx4��q��>���3v��I ��6�O�&�c1�D���,U��?}�����\��DŃ��	!��Bj!~y%��W�l}���ں|#(q;�_�#<@�ŌĨ�,fV1K�0�}lCx���	A��bL�!;2o[�lI3�*^_��,��]����~�>�7�Z��AN����ڰ�G��i�sY*J�e�R�T�J���X*�FE���!� 2��aZ	gQٶG�aR����R�%z��w'���2�K܀�E�=C[�	����Sdp��1d.�5�F���hn�U~�f\`�c��Ͼ�������ԡ���ӂ0���g�Q���7M� ʹn��1)�>4�`P��0�rq�8E�����\vf����z�)���?u�𣙆Ӎ����d�B"Z����8��4��$������W����D������ۼ�Gk�g��ݿ-c��$Q�K��O���aq9��o���p4��`�����`�Ȇ^h�[.exrn��a+�`�=�Ɣ�}�/VxI�� �N���O�����s�����xF�U�bFhH����6Tf�q�T�gIy/�x���t�O�*wd�Bu`�(y�R£�lӆ�k��ٽ�0Z׆>=�v<���~��I.�{򍧛e��׺��n�NY���U�`\X�kb�*ի��H�t΢�=��C�h٠Kk躱���B<7BN���/�Nୡx �2�����d�qH2'��]���˔�ã4r �.��y [}?���keEr�&�E�A�^�y��t���m�3���M��o�z6PR����/k#x#��_��pѕ�J�'ꑞy6g���N��MFKB�~2_�gL�A��!�2�e�v��zN ut\�AJ{�u&O��!�Ly�/J]3	D�2o�cZ�x녃KU��vE����)����c���T�,AO���o���՝Ǵ�>��R#k�X/͕�$C�'Pto���S��6�t1G��cf����w��q��6l���7Ҋ�MsV #u��ч��7�X��ʝ�¶+�F�Ř�*
����2'��Ŏ�e�؈]%�^��;��S�>I7�E��S�I��/�3� au����b}p"[�T��S��ʧ�w#�\�1[P���*؉'�ě��6n����Fa2@E����|L��H���*���`煙J]����:�p-:��G��0l����4����Z���jC��䪅/Nrh�����"����!�`˱�G�@X�E�奒w����H9!��,%�}nv��[:6[)BZ�A���|ɒ�2F�*u�]Sk�+$am�ۏd�j� ���e9gaӢ����
�qX� o(Q�� �b�廖:sL���4��3�P����E�cz(�T+{#a�:!�Ӛt���~h�ߓ��,g�eS���G�}c�y�F����K��(׌�F5XFS���m  !���r).?�ߐ]/��ϪYs���{�)��ۺ���(ٵ^���˛��gIH`�%�͉��+|+�m&P�$U���MD-�	{E=�n�����j0�$9M����!K�X�����}~��R�����N��Ҏ zڽ1�"*�4_�T귟�E�#"_��^��@I������Kϱ	S4�;��ܚ}AT��sSo�)+��d���r�0�����K�5����;�_���%�9�#k�i'9ܝ�of�rN���
e�9�)��q�n�V:���M!���=�{��A���`����uyT��&�Qq�����Êƭ@ߔ�6��=nΟmP�|i��Mt��L����v�>���p�/w�#��A'�(2:�l��1�A�#kÓ�B�~@��o����G��m��Û�r�+����	T����w�1��@��kê�IJ�a{�}�����;�!��3����k
�f�4Y�Ӥs�h��s���#r�Pm�S�mAL�Z0O���.��y�`Z���#	�}-���,�µ���X�8�d���y�*98*��e��Ќ�d/Ahz�?}<�,C�����#.V���x�[]×Y5L�c�N�����DD�0���˼D���WA�E��C0��=�WP�V R�W�cL����VUW#Ā�@�amw�Vv�"Ǚ
��AQ���7%3��]�Q�+폹��(~P�$�4��\s!�|N0!=VYBm@�eK��ʣ��{D+ �L`�{՗�(t_t����iUC�&��/��G��2��_�b��Q�Ȁ7�G��$���E��_�i�Y� �1M���GSR��H��pz��^�q�n#ugߕs�*Mf3��є�'{3�����(+��i�������\n��nv�SP��r�Dr��.��C���պ;RfI��=ck$p��o|r4��Ou��>�g�e��IAņʞx�˱P������O্��-�c�&�o���?��'U�"���0��T�&�G�cI(��U�d�%��74j*��u�g��(%��;�J��97����<h&y����h\7�k7��O���~'tڎp�{��%�:	c�j��Ƿ�f�]NOW;�[�t��ڬ��Qj�-�Ep{��cA;�����i��9���	/S��:\�!Ռjo��*��[��ǕN��SH�N۫dw��&�!��gW��yp%�J�����Dp(MjAVmU����\.�}*�4�J���!����6���S�	�PA�V�!�(R�ڌ�q���ĶJ�y���Ui ����o:⨳4
'W�v!��ss%�o=������8���.��!d~�F��Q6�݌b\�,�ɉ���d`K�Ŧ��A�H&�>T�����Z�W,=�ظ��dNޕ����P��!j�x;J��p�	��d�,'s[�3�6'��Ko#ȗ�s�n�ye5�u��/����'�����
K����X1ή�0+��Z\���SU�i�r���~+���+jF��>H��gP������(�� �K�`^�0���>� �Kbm�]��:T/��b�\^�*�]�A�&�h�b��#/@�j��s9a�;�/����0��� �l=�%p�q�@�76�p���i�G���8��Z���|:kLI�ּ��q؉��B���;M
[W���,��
�T>Xa���{^i�u��H����V)W�w�3��c�<.#g�p�a��a��	DJ��3�Ӊ��.e`�Զ �A��|p��#���m�՟xvI�����ђ������?������[�)��B�_�߼tO��I3�N�-���;���yˤv�E�>'��v� |�Kiz�z�aW�OF\���K䮤���>6��9��rb�־V���a�!�B������Q�VI�����9�ٿ�
�o���g�Z���,C�"rz�08A
��{v��g{�I����'�M����5������j_�&v}̭�֓j�].�We++��]�| ���5���ʄ_�qb�����O�%�y�7ԹU�6R~:�-
h�50�u�+��h!�<�k�듎��Bma��S(�y�Q���$L<!�	7����d�x���!�H���3Np|̳�(������xA�c^�q���-�ℜ-�d�y#�����Ih�Et	iū��i�6���`=4�R��o*w�)�]�fxY7l W�*&<:V�	 -���5�J%�8�W��.�s��B.�q��W�Vj��v ��I;�8n��ѣ_fo\h+�~��jk4�Fla�<�]����I�\�E��5�e*=��K�'�;kVA?օ=�c��hYv��is|'TV_�(��Ze��5��+�S	�Q��j����ɯ�s2�����y<��c�Jm5��l��¸R�wMI�n��>�^M��x��N9*?��0��>��"h��H���K�P�-f*�hrx��k����,7���!U��GT���y����T�1&o�}hק,ҋ�L�_؇��Kߥru۬Z@������ZDl�s>S���g�+�(ܱ���:
=J�x��pDVW��&�E��;U"�dO��\�e$7Q�YC��qk,:�r�p�R�ϑ���*���5�����:���������M5�1��Q��$MYc�m�����	���!#w���K
m|��$�6x��(��˃?��=]Z�}�ԗC�x�&����-P��������F��DC40Y��f}��^A�,|��9���u�_�s�2^~;t�Jyn�����:6v1�\&��tp���b)�g���*9�*\زy[7���6L�"#�S0��T�~�@"���P
��jw���s��	B�`7dneP���;�gH��f�,3v��F?gᛡ�k�;�M\1�f��]zI�?�W~��ǎ�NTC�l����%��.�W^��Y���g "�{��SP�~�I�P��B�i�^$�w�6�����u�E��~Ӎ� ����FW�S7��u��1�:Uqh�����z�+��=�,�z넀:g�����B1�dT��9��=%�Kq	�����x�^
��j��~O�x\��o;�����w,�t0�
�|��Ev��z�,�n~.`����$~ޓd�#��+E�����������)�0���s�\H��0J�<"�������P�4��0Eh��xL��Fk�Ơ���/gŽ���:^��!��L8�`:!�Xt��|})���[��Ҩ��W'���-8�O5`��z��Z��t����pb6�kk�K5��Z�K��>4'�d�Ń�k��f�gy76%m���R[�%;�CW�]��\�0�_��3�����na�|$\<��l�s�T�WCz��?�K�-{-��,�����cWu��tC/-�g͟ԭ'@5��3[5� _�虩O�NC�1ќ���s�t
��v%.V�0kc����뛉$ 1uG��.î{X�1w�^��ڮ_�^/ߝ�4�	��P�	��Ϡr�,T�!�tT�*����,|����_MB�v��������0��C*g���3R|�?I��A���Q�B�<T�E��SD>���&I��\cXL2�+A ��9:�J\�����1Nj��M}�}�"p�B�F̔a��L�"�B$*���:�K�jfX-�Om����@��\)$�N�W/��!vc�ywq[j/A�Ǡ��|��b�a��L��S��@-�ZMw�t�9vʜ�Jx�`r�ӸP�O�)�B��~�Tް��UV;�%G˲�5>/԰,J7�/
���ʧ�y�>c�k^mԎ�Pn��*W�ޢ��%oﴌ'j0�� ����E�K�B3
JC9I�$����`���"8�h���k#�3�q�~k_���������f��
�9o�*]���F�M~J�l���ېI��_D�t�~#K9o����o�C.���e��$�����F�z��4D>���7Km��v�J�(�Z��Y8A��V��愠-7�Ϳ�'J,R:()tk"�s�<�:@;�)��tH{�_RR�-�?2d���8��m����+yޓ;A�R�ַ�?�S�����>�̄��e���)�i�&������ʒo����JX�:I�3�7`�$Bq�$�z��j}IR��Y����묰�m$�r��ꨞ�+i;�P����=4\��_В�Ϥӛ//�ns��0�[��s���h��D��Oa����Q��Hdh��)��׌����q4�,���R��v%�<�4�%̓ƜCUYh'�E�|=�@�]��h�Ɣ(6*�u�g��.|�N�3šR5%񔺣��cA��.X'[�8�#>����ᓭ}���dP�ǫ@*�k���I=���`|�}�%�l�~���E<�Z�"U�O"���ueڣ(w���jd��@M�p�E��κ\�+h�Y�(����hxO8�fU&B�N�}���G[~gv�^r ��I)�ɇ�0�� ���Z%E���Nm��ɸ����n��6�q�[M�u�AD���V� �)�?ߍ����#a$���7� ̪����n�ҽኊ��d[,�)E���|2$\���*�5#󸓲*��3yo!0���k�Imxf�zC�R&�yL�x@8���3 ы\��N��D��Ҭ��Wd�|����1}��u�m��w����##{WC��V��6���N՘�>D�r�(S䱒�51�s.��r���1s"���
5DY�N���6D��&�`,�F�'��d'�t��f����fP���b��X�#�z���_��LR��"�t�|�Ò��.w
q�Z���~�o�&�����b���б�"�?��}�+�Upx�N�������ANc��n9wW»�f�^�LV��.AC�ګCg_���V��g;t(�VL4tS�ɑ�x�;��I�P �_ "���$x6bz�!\��6��$ ��Ȟ��P{q\����(��21K��ɝv��!_���*_r�i�����.ȑ�a�R�f��̦�{M�k& �������8�$�$�l�a��<��8'�;�S���U���4�_3B��u�)u�wy��#2���5�h�W�V�+yc"��)����<T�r�ԔQ��y�����������,���H�6�+1�&m\� ��P�����0]����,��X(�%?Hg��靑�������e�L��2d�X�P��>guvS*)���0O�<�
�j���e�����S��S�m�}�y���i�&I��g��^3u�N�����B��옛&k�}�pԚ.� ���[=g��;&�2�C����T�)��P�ᒔ�V��>��v��q�H9�]�pJ�+���*������rT*�����b�81�dr,�/a��x�
!9�s�g*�	�!��R\f�*��J<�R����Y4�;{���B��;���'�ȟ*�IIc�vc��m�[�W�G��K�F�,�{�h)�8�����|B���c9���]�ĊF~ŕ��k��0$UP�w�|t�H�xb	i&<�cʽ.l��z-��]�MlAbW���p��4D. QK�OzX�}+���z1nD��sD&V ͯO�����`���dvVf���:���
&����/�>8��F}��U���/�E7e�ŉ�o>PLT&�R�n�Ł@�Jϣ|Y���2h�#�����5P��d����E�Đ� )��
$���T�lq���|�V�9#�U��� 틲E���HH3��V>d;�J��8ii���z����gN,�a֛�X��	TC12Km@���L�K���w��39�}���-�ȥX7��~���U@<�bc�݂|�&++R	>���>(��)���+���V��9y_�zK�'��`$�@����d	����kG�lu�m�Q-0�����@�Rcm'�����x��ʐRΕF��N�ʴ�2O?�C�XV�Ȟc� ��<����.��t�C��`,v�{�E�8���>�X�~[� �㐖���%rU�A��h>�g\f��kP��j̍j|R)Jv� l���d�>�S�D=�q/�9�a�Գ�N�^�Q-��|u�|(:#چ��E������
��z?��d*�vY���o��SZ��~��������u�~GL�t~��I)��BOŸᩜ�׉A���O��i�ϖ�>�7��Vla�x����c~5� �a�3k�Lk�s�Aʩ4�z�a+����<�r��Cl*>h��)��C]�M���r�U�:�z��"�N�	�"_~F�H���y���t\Mi�C���
i���ȸ %F� ���d�e�ĳ&N�I����4vJj���*����n��BǴ��ւբ�&���oC�4���%��V,�1�-��<�ڍٙC���o���O(r�ƪ+<Uܩa�����U��>_I��rR^g��4�z�e�)#ɶ��Z��.y=°�p$<F�Z_�u}���Y���S�A�H� -�4��dCP$p�a0�VZ���#������N ������\�cy��R��f��I()<��^�,�&�Z���x9��\v�R�<3sv�+����T�,./��D�bN��꺺޷Ӛ��p����D�D'���B���a[��@����4�q�Tb�6�΀�� �1^K��$k[�[Zm�n�ϟ���!�i-� �ۄ�&t�{���u�w�L�|��'�ro`�8��[�,c(*Bb��0 el10J�Ӣ�~kQn�L~�~���i�8  cD��֨�<����MJ���:\���^?j�;d��HO��v��2s1$x���O���伋���Q�΃[�7N�6"��F���3�VfgLt�N6d�8`�w�μ�w2Tl���8A�ܹ�h)���ƚ\�\��@��8�J�x�@��4�Z3�<�3x93=m��{h�Y�L�ͫK�O� �f�<�����ό��90v'Qr2��g��S}.��a��Қ��W7�J�6�k����{�SF��/g'�����˼�.�����hv'?�2*v�`���<�&�4T�fg��#0��g�p���R�?�����ȘwNQ}j8T�[�U��̯���b;|٠��q0:ٯ)�y�Q��$4$50��Z��gB�p���Pq#G/z`#ᴶ�m7�b�q��&hw��VJ�_����/ ���X_y�Q�� O�np��l�ޭMw��ъ]/�Nb��h_
�Ah�WX�"{5;��CZ#ίª�dj%��jZ{Ŷ��OJC�+�H�J�2l����Q�����a������|2j4j+p?L��\U�8�W��v��9�`�#�#<+���q���ry�;T=X���ܘ6�7��㙪��Pi�4 W^9��O��΅�IJ�G(;h�Q������QnGӴ ��[>%5�w#wb\]P�5�KP��3n���������f.����_d�uw]��5\��)��������#�dn/} �̿/R㔠�	C�@�� ��r�sZ����N?u��'����@`fx���4��.w���P2X|#y[^�3�
�D���� � �4�4�$�s��Z�&��\���f�E+2☎��QΠ�O6�פ�n`�Y��Em��5��]a�����@����@R�vu� GPٮL��TMh��nv���̒���Ȍ�PWئ�U*_Ϭ#�\���QƊK�(o��(l�a��߀�� �|�V�$���~[;۴��_d@�luޡ��@#�X��������Sץ5�Xz�-K�8�X��Vy��û�]�-I��K��X'����Q���!<�G�H��ԓ���<y6�W�^7��e�l/�ra��q�����n:ɞ�|k1�7���b�%�0�����B�P����bׂNO�k�Z�yAC$Y� +�JI��0�����y�[�����`��6����tM��C�j�|�+5)��rE�a���Ca:�y����E�Q#�+j~���l���|��M\�7w������hH~VZ{'���9�|�z���B\?�foE<�G-k)!R���pxJ��1��P�%חeM�= %Ų"�	ӣ�����/:��<5�py'�b�t;����fe1A���9�n� �5�z���ܢ�W��
�Sf{�@��O��7 V�ѿO|6�P��� �O&7��b��I��K�y!4F8 �}y�W��(8���X�TG����ݯ�O��� �J�Շ��}�*a�<�j��I���D	�CQ��d��OԚ�Z�[�͔ �։h� �P�bdBt"����e/+�G�vL1#�˅\�ڮR���e����>ɢx\�}�����ȯ�QR��M�F�3w��[�Lau��=T	�N_�z�q���a��^�e�[Gi��@��I�*�*��P+��ZБ5��pH�װz���S� �7�P������}�����6h���I�c�C���?VE����6��X�[ލ�	��'G�Q�_׈�0����\�1%,U�߿]�g��ԜF�<��C�TtE�27l����L^�,Lb�q\6S����N��3Ю����x����A�BԚ���r�Fm�lށ�K��O։�X�G<�V&�+�O�u�>h���x�Q�d�ǌf˙��Gr�up��&����GS�f;��Lu�3ur�Y[+�=���D��ٻ�N��� ��O�@6$A�Vob�G�1ۅ��ZA�����'�������?~�d.10��
۔���H �uo�+W�QJ"Z�V>s:�C���M�-��
J�R�d&��.h����X	O�W!VB5���`�7����S�D�d
(`p�|*�ٹն����� D	s��w��y�ƺvd�Ɉ�ُ<|��'\G`�Ĥ��j����z�Y.���j��M�|b�l�赯��\�1��i��׮@����۩�����i�kE
���(kp�6�a�5"ลK(�Ϗ�d��ep/���1r�2Z���2<����������f�'L��!��k��?fJbћ�8��������U��Uh*py��N�VVh�Y�d�xgw�Z��U���6s�	�3��]�,j������W�UA��}��4LB>�	ߧ�����d8E����~]ɧ��NJl`i��5��g��ƥ�z<╨HRZ]�H��ݒ�b���i�yHo�'�'�GW�n��H�XY)���k�D���Lbd��c �U�g��,���(^r�mX��j�~x(���ۆ �!m�1?�L���#�p^M��L�\*���1Q�x�= ��~�ϼY�K0�K��ڷ����^��S���XJ��eЈc}�s�-U�`9v:;@�����ԏĞ�����5�� K��{hB���M�Eڙ�����g�x�3~|t\8ͬ�Ğ�%�OC�0TGO��%OC��/��<�|�Y�(	�BUتA���ݰ��G��U3u����n�&���8DI�1h7�г��mE
e �pr�^�#�$b(Mɿ���%��^#�*Jh�r�^ۘ-�^��-��G�Ý���>�^��`Z������-���Q��h�s}$������"|��usKb_��1e�g�� WΖ��<ت��'|�ʅ��t�0��%��La�b7�p���?"iy66�����N�~��wLҰC��]z��`�xH��,�sW��DU R�A����?dӈ5���aʬ�E��n>�T7�x�^�%��g�����4Di6�9��tIU2��pdFԧ��#�R	)o���P��eG��NБ4�(�����f�L��)�a��>�Q�7�Ӱghx'��0��N�y#��Յ�M�rj�m��TU�ʩ�=��^[�����R�@{.���r#ydX[+!��F�M���N�kZ�P�Ȇ��V(QB<K�x�t��c�C�:[\ŉ�L:��?҂��� ;��Q!�вx�芮���.:�<�0=|l5P[R
L&56�sy`�/��p��c�U���=�1Ȉp��n�e9h� #z $  ���M���?�/�^���X���r���˗^o���;/a$��-N�//��u��>���YsR�n��ߜh)b)�q���*�������͛�ƿE)�iZd�#0/d2���&rH"���I�RR�X�e;��9��dl~j�&�������T
�s��Xu������&}Q8>=��LY�ЦB���w��(�m�e�Ӈ��������kW�L)��+��)�Z6l��:yՙ9�8];O����IX�
��يs~�ԫ“БR̷���m[���Tt>w�F�P������;���s��m�
���<�vñ��5oJ�|�0׼��啺gRr7�B��Bc�>b�`��x��L����D��
v�T�)��	�E������v��ǎ"B�~@�M�ŝ�[j=�I�7���b����t�Q�k���.,�*�u�ca���v�u�sk� �M[bf�� N_
�gJ�H�f�pe9Qs���|
�a�8२4��-�7v�1$oB�_^�@��k�w8����ǈlҋ�W�t�Du��U��A5���Mk�����?K�rL�6w*�sb�Փ�����%�F/���"t�l���|&�n{?�v�9{F��;%w�3(��D�QH��`�	�}���C�IM�A�?�m��l Q��O22��4��p!�x�t����M��vH ��u�(]���J�g��ۼ^ �T2�ȕ����%�iȼ;Ti'�@��)����;�;�L7�ITq��)���,�N����⤘xG
9��}�3�v�D��H����2�-�AS\��(!��@W��WD�����N=� 9ʇ�Ⱦ���=c"����?u�h��P�M�U4�Vn�� Qԙ�E/]���ų��\��E���lM�Q�mR���9��L ���܋"��JvCs�S9
�v��:3��������մ�A5�~^y�\���6�OZ�i߫�N�� #`�I����N�gLqL�6_��vЀ>��Q�E*�q�W�cCa��x�����_�|��u�*�O����ri� ��\
�9��ú/�ՠ㈋���D�(��ާ�J|�w�U;�%,��/��_̫%V�!�<��"{�������F�\w�y�ȡF�}<�����<���=���C�X쐽�!�˛����gx��-�ʔ(�Wޭ��a6
�1��ӿ� *,г)��nȓ�B�j/0`+��=�0��GZl��e��<�uPcg�*JfHE4q&��E7�����~w��Q�o[&R�o��ၻ�K�#sɊ��حHM���f���1�����Ő���6�Go����ga�T�
����՝S�̶�?����.[2i%����T�Ig���'�� r>���EFv����_{�L�tu>��/���.{;�9 # 9�~q��W�ŉa���9��m�B`9�r{.��&��]�}	���?�XO�y��Y�%�m�h�ް�{O_Λ$��Dq9�y(^b����O��1��\v�xV�Yw�>Oĝ���Z���o�Y -�G� H7�D����M�d>��RhS`		��-�u����7��]��Ļ&5��+	>�g᭤��`�����,L����OFL#[��#0�j�6��[���S҈GO�No������Mo��"}�<� �!EĤ�"�1�w�78� 8_�Y&����X���U9׭�I�w-�������R� ���'D~��Z�M
Uq��c�c2��zsB���e�|�2$�*�,Ф�ٍW҉��4\�wsN���D�2�]��M���$��V}��S
9�Y�%5ϳr���9䱞�.�tļ$o[)�a#��)�hp	*9�M�#@ay6�:��k���F��jW9<@��
�V��{�F6"U�|s�`�9�d�5�1�4�zQ�:���q<�[1$_ݔ�:S�M��`
�w�9�O���&��y���x�SPx}Tn�'�oUrL�.�9l����9��,ӥh�w��4-a��/�?D��J@Lep���W�1VL0�<_n �)C�f�@PϽ���v�7��{zR�R!���	9�%�\�-�_@�?���[ۖ+�bd�IC���,⡪l!��?����UB%��גּO/���k����٭(T��#'TWkP�޿�<	��_�",h`�T�3�,fkN�;���2�T�@�C�Z?cGTjO�>�'QuǶ�Ta�/�
���.* F�}��'�~K�B�c��.���c+���umR��U�O:'pu'��=N �"jը��(��T�*��[������sE>S�)��Γ���ݨA�P�U�'������l��+uV�`��4I��'�v�e�u�XlO��Ζy"��+3��P�d��<���.,k�ؽ9?>"�����XF��?\ˈ�|�9��;�hr#���f,<B��$]�C!h��bոo@�{ײ/82�rj�D�=�:2���I$�+v�ܙ�	��\۔A8f;�X��ә�H�~��iSDi�X���e��ٵ	�g��R��&�ɺ"�]��f����a道����Vc��xg$�.�,��.z������K��B�>�#l�5BF�d����LX2arQ��ѡ��=�?T�t�,��I�UO�Ҿ�)MI���Y�Tm@�q`�ZEP��pA���g�ɜ%1����l���y}ox�چ\�"G�/�s�l�y�8E'^��RU
_��geٔ3�Rv}�f*0a	I9�.��dˍ�.3Pb�k\f��37 ��X������z����a�Np6�O�<�\$7e�0R$
�I Q���w��0�ϛ	���P&�cj�K�����3.��MMؑ��a������
!c���C��z�D�͞���]���?�cAvz�0m���\��mm=��&�яY�q����|çՄ��4*��WD?@��|g��J|�e�9�Pe�A+74)�4���3>��� Z�G;�|�h!K��G��(�Gl����JЋ���qjOh��iL0*v�F�].�h�ᠧ�)z\�����]�����n��HJ؍��3F[G)}�s�y0zu��u�����͂s�R_ն`Dg�x|V��_LC��m��ץ�����C��~܋fNZ^T&^ԝ`� ���T�l���,"� g+��&݊��:
�a�)�\�O-ȓ�Y��o��J���vϨ(�QYqW�_�sO�6�J��f8Z�x	)r��+�)�Hc�J8�����p�������+���s@[F*v�z���ᄝ�{�㢣�3AYP�z}��mFࢨ���(�"\"z/��4@�o�7������6��$.ˉ�G��	 ؐ�i�Bd�c��qx�D��]��V}3�R�Ul$pw ��.#Z��!֚J�.g�����l�\�qz�T����f���,�].�(D�¬Q,�����"A�.S^fF���{qnט(�%�m�$�T�>,i���B����N��FH���:��lu�>~A�����|"|�:�ע��&���v�ͮ���?���dQ��D���t�+�d�1��8�\��>@ω��]k�m���q�K*��"�=�)�M Z�c����>�P~i�C먯ޫ����|x��t�ж��t8��3@�o��	����|�� #,~:�?]�Fݙb�S,��$���T~P��7��I����ة��=Hd�n_�=��E~�n�u|�N��������X*bY-m"�'�����z��%)�M
�랥hމy���0aM l6��e���i*�9+ߨ�>=Q�G�<���v��ɜ����+�ѸϮ��U�OH��[�����B�6,A����t�,��#�YM��\�b���?n����bk�jI�T�l]�5"s�p�BI#fТ�h�PR���@=P�Ա����dL�xx�-���y�>q�7�}?/O�ٜxB�\1w�U�=�	�Ŧ�Y���:��<˯���N���X�W�3^�{� ��/� �j��XG	�L��M��]3~B`��򾥲��v����(�s-���Zgy���%:-���M�5����b���@�_�C'cO����&{G���}!c�k�_���7��:���;�9�,��0�\Vf�� 9��㷫��O��`q�2VU�����N(sO'������pC�q1�A,=v�(�"�L"�{�ȃ��:��C�P�0�t�5i�@��n3.���""{Sn*���$���K�tl�K�!��X�.]����{)),����9��b�D�-�|j�[��5G��΅�=�Ҭ[�I���M��>2RK��)�_��j�=+�F29��Uy����#�����l�Z��D������ǈ&G�
�4�P^-��_"j�R�٨@?:���/w���B9�'��.��K��}��QD���wk�ׅu�Sv��K��(�%��Ca:'�_�1ʆպj�[p-S��)^s�$͚�E��D���)<8�tA?%eaz�@^����n�ҙ� ����TU����w4E\��Tg������r�N����'��kh&�P�ߓ.W�WeD��kU�/���)E#|�/�t����Ԩu�b%��X4�S����M��a00w��TQH���d&��K�P ,A�7���6b۳!AYXO�*�!��a*�6��w�["�/t#��(�>���>^���V�^d $<�{:>ܫ��sRF|�uh��"F�6�dn8�T�V<�.m7=6B�ά��?��O!Y���D��E�)HRk�E��	��^�-�U��1*��b�$��ށW(��'�*XNӃ�ܟ���Ӑ��&[��(���s����%OۦaET��� �S��8�i���~�t�H�c��.,�(?���1 �0�1�6���(��s;��7~��4
�V�0	��u=�K�j%!S�D��C�v��
�K��Td/�%�!����r����Ø�8��RXG|�ϐ�Z v%�WO�?�9 �0�����
8�L��
�(�Ä�Ń˦Py�w6�I�l�)�<�`a�~(t�j�+�ǉw4��D�H80������,�e��;���.�#��V��������aK��/$�~��&H��*��\��n'b.�2�d�AM~s�⬱��M�QOAY����ށ��UF=�)v!��?vI~w��I��$g[O�e�=��EP��U(�v6�sHU���v�?��� ��J�:},t��S�	R����J�>S��)%����v��l�K\�4`���ӽN�ۊ�H����Ū(T�N�z/�!�*���i��KA��nD��������H� Nb�A^s!�֨>s�&`���������R�����Ji��(Lfeb�-�%~d@r�� �e����A"�,I�=��lʲ�b#�g�˦t�uhU˱�;ǟ�]4�ؓ�GS����vR>b��:���d���$ǠN-[����.=�3�]�����8C<���N`%�~a���C�<ҋ�t2����ٖN*��¶�UT+��f�|�o�~���O�:��z���e'.8D�-M E�1��O��f�[�!���X�3�l�&�ȳ�x2B��3!STDcM�\�]%�A����D�o��@|zqg�Ɖ��`��pa��32������{@l�B��W��Ci.��-�;$����
V����T`�k:�[�9�~t�6"ἧ�~����Z<��2v�鬃Q"A�)
��>/�8C�]�j!�a.l�1�"맕�1�^�1���]ßq]y���3P�\�y������q�L��e��م���-��)����A��Eue�3gA�}l�����	x��G�~�՘�ʂ�m ����/$O?�� ɷzuO����Ipq@X�Mg���>͏H��s�o=@IY��U��"�@
�e������Y�V�ӝK��I�|z�φs�o]��j(FP4��+-�f��H[�{-tI�h�%01
Tێ�ؔ�iď��X�)
2
�f��nQ8d�c����.y���<T�k^%��V�����<�a�v��d�
�t�F��:JNW4f6�ǘg\{@A�j��[`�Aڰ�$�Ա\��!fdU%H7�Mkx$��o`��rݹ`)]�jı����2sm��f�!A'Ji��9�z6����z����6,/x��}2���3./�c[8(���� �-!Im�06�+�RC`+ Ϋf�j!��,��b"w�����L�?(��$��B��9\�i��`�BlWWa��"o�@B�˔Wd� �C((ԍ3w���@,��fOlO����h(�/f5���{V\�G����-W��F�N�^�Ut�_OV/�Ή�[�me
�Lv��2����K�8G�y@�k]f�yU�y-�2$��i�U_��{2#�9z�ONĤ�Irx��"��d|��5A��BƮ��i4*S�&���^�p��I��پg�����ۡU���p��T�]Bo����xCt�lɳ�ZV �C��Rv?��þ�Q>�NN0A�}���9b�΋��z&U��r�7�
�s����eػ)��BK�JF�Ts����G �1���`��z���5�+�")���??��]��M�a���&ND�2�\�;\�I0�G|�����)G�U�e	��G�/��8I�f�_s�~��
w�ջ�mI�aCb�x[�"��y�"�m��3>h���G7(��I�9�5�t��|�!����b?3S���h��	�
:��<��9�Ҿ���Y8VI�=}��5�zdI���_�!����ejNM�H�c����K��C�:����g�W* �[H�Wx(/�oTqV��J�XS0��[_+���PS��� �|�L�oR�t�;���T���Ӗ!���hk�	8��P�6���U�,��D�i�/�A�v�ϛ�[k���h7i;�����ذ;�D��L����aï�1͢>�+p�����,&�;�T��\>S�?�e��yL�.�Є�Cޚ~;�_%������ec�����n9��Y�ˎ�T^t�c���Te�R-ȟ�ʃ�^�:�Xcd�S^�ы�B�J*��?�aBfxZ;�K���g���ǦS$=kN�
W�
��Uyn.�Λ��˨������˙�ĨU{�a���r�H��������5k�Sм��.TYe��ކٴ�!MF�h��=���%�
�����荿=2�<�-cn���ALLO6WpkTxMO�ࡍJY����!.�V�1m��w�5F	���L)m��ꏧ�zcF���������N2s�z�s���6��&�7��H�KQ�)D:$eL#)����y��?�����Ꮟ�66�)S���d�bZkfة�h-[T��}#���������]�?��5I0p�}��?���q ^��Fj����D���0�
5^̋/����D�A��׷��7�Xv���|6E��rU���ȞA}�ޢv�ɵ9P~,<$1�7vm�Q&9<9��Q����uu{
���qÊ��X.y�N𔑘�W��j#(C`&>ED��D���t�Xp�3�+Mo���x���:2���m��Il��=Dl�#�;�ŢL$�F8¾�1\k�oLm�!ԗc7��F+����\A�J�P�m�d\4��������.i�ϪW�x�3��/[�����?��k?�7�uKS��0=a��s5�(F�֛.�քIb�CR�3��ӥ6s�Y����v�5X�0���9݈�C�G����Jk�.s`���wo������ ��ֱB.#5��a~O߇+��X����]����Y�E�zM!��ڨ�h��s����;�@{�ПAE�Ab�C�b	}�}?Id�I��Z"\�6��#7��7�
\@����`�d�cz�%\�;�?�w�8a>�9޹:UF�s����K@��H����x�w��S�%	��1�(/���r��c��*	���-a$�s�k��PQ�dw}P!	�w�tV�=�������-8!�K�5u�@S���ǡ�8iW���N�ޔ��uDN�����Ar6dܼ!m�N)���[b8�����Y�Vߦ�	�����K�H��mgtiC���>��hB��Z�n�웝��T7:�^a�Bzc�L�C4ь�%��y+�"?t���Y����x��$O��5ɉ�Pe�ڲZ<3 vL���lH�
/X�x�;3�RSϴʛ���peqTd���nz=]YV؈�B!K�㾆��/� �T�u�#Dxyq򩮴O+Q��c$�^�l!K,�1�ឆ(3�T�/�z�wc�Sɍ���l�����f�o�ឞV��&֥�ɍIl1���z/�}`�\걬����(|'���l����T;��5[BH\��Zy����?���aE�%��A8߽�ݓ���� �XHC���P�9+BkF`�GJ�O��c���+��.Q�OZ�f�3��d�ߩ�����V�0���X��Ncc���xR���&�s��\2⁂�M���i�\)��Ә�[Z]�N ���f ��0���i���v�j$Y��M�vg(34*RY��E7�(`H0���r7�J����Uc��@�f ఁp<I@J����c~&":�Z� ���\����=1^�GneR��t==� Up��$�[��MѠ�A��a���[u�)�E�W��w���'oy�38�eD�Fk��A �AhJ3.g@���.��^'�(��u1�5�v	L���l�"�a�ڰ{Y��y��l�$^�|Qo�f2�Ec��3<��29PY�4kR��D�O��?�sG��go��$�J^���0,Ԏ]��w>;���9�A�d�ڏ�nwɡ�RS��+�ī����Lf���+P��ɨp��������y�v��b�öb�5ˋL��9�%e��d2�-���C��B�_�����H�g1q�)��ߛF���(�ƣt�=�Y��?���:62X���/����n0��@nҞ͚XB��F��
!�z hFK�40JTqt����ݳi�S6)ka�ϝk��ՅwFr�l���F�	j[��(�y�������-5^��3�{ip�*�.-Q�lʥ�-��`!�b���W)TC����%;�A[�#(���OЩ4^����JNQ�S����̲Ė�ܲ����q�����A��i�T� ^WT�t��%�_�)�q�~�N���  ��
�$2��H���'΍VJ�|����������:�SH�G�C$��=�Sv�8|7,���� �j ��&>)��<6a®UUF�`�H�������(���][(���J�ģ�Q������2/��+ʰG��YD�T��#V�^S�ɻ��t����<����U���X�a3�<����8zG��r��Vaa�q��SZ�^g��y���8ku�����D暟~�����Ԏ�`<H����+����6��8@�Ң* 7 �s�����)�'m�(�+��w��t�^0(��$��a<� �����l@~�Zy���'�:Zs۟#(mLM	�My+��y1��=e�?����� �R��/��2�O���*.as8|������b 董/r԰��o�
���{lD/p����O�/����*�n���"�b�V��jΑu�<7���ؗգ�k��8^]㿒$b�x�_Aa������!�)�K���A5N���Q8M������3�i�3��fD�P�z�Yl[��O8�<'I¯�9�m���4fR�J��{���iR��udgxu�M����G������=�HG
W0����n7Ɣ���C��;�]��t�1W��q��.+-��` P�n�	t�(5=�A.*��X_�o�ֹkD��䩉��8.���`+��~��ʹ�IF�L����2�K��ߚ�H}5���?&l���|��D��6Pj���ب����Uo��U�w�.=FD�5�$$+|��Ȣ��i���.�����F�%׫7\w�,��g�E�p��������VۀzM+�S�$	X62Y��w�b`�����`�A���S�7�U�2��<$�/�}\O��/��Y�Z�ã��C8,n��jN���F�O�R�<c0= ��D(X��fVԤ���xW����xk�5L��4'��~{��۞�e�c��NT������:�y�0d���v��=�-|�#t=��:X(���l�,0�V��u��*��6`HM+)�[G�S��y���|�F��)I��d���2�	��� �P"b�t0`�q,�P�	���uD34;hB
�i�3�@�> �����O�ˠ�l�����"/�����|�f�)�6L;�%kLSo�����me=�&M�Ɛۚ5�L�7u�
�� K��]�h��{Zs*�RW�)tu2Q�<�ls��v5L�v�Q[�~�~64�K@�rqr+�UW���kQf:.���N؇�\l���lyF,"BB0�,� a!�:w��S!(�#sv�_���<�~������U�+�<�.�{����.��53��Y>�5��b�[$m^���) ��itA��G�u����T8
1�G�y�,/M�)@4�4A�i��)��52uP�0h�T �	91w)Tt���+����w!��G�o���0�ʇ;Z!lQE��C�_@�2�����Z����:���@hO���k��W�Z�jFV+}[;��Rz���{�J�rU������e�R$?I	F[w���:�x��+�ݤ<��qm�0�9�,g�SE�����{�6��s��0d�����蠞Q.L�k��A	8����@�1C�8oEf���a��n��W�Gk��C��ܠM,�u�?����H�TRr2���Y��F��|������v(d�}�~�⵮y&�Rƙ���%���5Ɗ���5;�P7R8�4v|gm�+�.
��"�Y{�ya�8��p���sǒ���/Ę/X{n��*�2w��Ӊ�w��/@c|pӶ��$�mr[�Ӄ�&����D�&a���r�)�o��S�S��#������
7%m����m/���;�0�FN�8��*�@�V'��ͦ�7�������	�)��o���m]��Frz�DBnK�P�_�R��5�0 �<t�n��:���^ޝ?^��r��mer-���bv�@F��\ߜ��3�5�2DnFe� �=���є,N�P��f���@|:�κN��E��L�����4�q5A�wL�j��F��,#�\V����ȧ9�t9 ��êv2Y󼕦몪�y����^�8T��o��Π�~�XC�l2����0d��3�;�k����-h)�Qަi�������d�s��Wo���i��\���y���!�S�S�PH�^�"�}��請|���$((����ʡz�
�v����z6�3D�����
�w�'�� �����H��� �|9��~����M:�����ӭ@�S��Vh�7����� �El�|ss9�s�_�.�U��Z{��ߚ�=���?����1d�H��i��/V=A`?v��_4��������*�,�=f��M�~]^
ꨉ��2�{x�sO�b��@'�8H�	�!B��0g��x��ҧ$��N�䙴lcBr�A��<Oۀj&�7�Ԟ[P�`胲O,ګ&�6V�[��� ��w~�I���D�q�ȉI�ٷ����m�=��$D^�k���8ې�������l��W{[ߒ���3ڡzOb��"�Z�
[�YS^&�G��l�+�Y�2�#KDy�/�?�'|d�䄰(	���~�\/�D(LHj���<�	a��Yѡ	lqhx���4]`C��'�u8��aX�ڠVn��=�o��`���oᅎx��JH����h�3-������=L�rI��k1C�!���mG�7�J=%߭�\�r�k�F�W�����&��z�Ջpi'�O�͝6�@�C���ٞ|��zŁ`2�6Kr��	�DzS�b��Bw��?��N2��NHՌ���[��k"��N��u���G��=]ED���yj�J&�9�X�CJ-��?�v�1'��oWZC<��-���Z�Ql��������?)�[� ������}�.��Z��n�[<��<D>�ȟ��<�ϔ _1�l,䶾�9A�k5�./�	3>c/)���s�(GΘ���F��q=�س%�U��9%���ބ�ʓ�5�t Ѿ2U�FVf�.����I�u�g���k@{��Ps"���c��l��i�(Y��ow�'k�%R�XTBڔ7���b�4t����P�{h#�1Z{,���&�MSI�ݧdLRw�V7���T '��2T.-�Fww`K$�ڨtS��m�LR<���u��zv�5��U��ɼB{�����rn��c|�� �|st.�Y"SΊL����7����TEx�����_P������솱CM��z�X�� �>�$�(?�����4���j��Ř��;�/q*@���Oe����%�_�B�.����>0P�`S�đp)E�H�"�3�$
��|L+2Z�4:�W�;�jޑ���r+��#����@�#��N��=��Sѝ�����1m�/�X����BJ�غ/T��lL㮧'
��t�bE%��-���j��?X>����n���zl�N��Ԡ�{�t`�|�"��rT:�Y+1�3��1�Uc
ƒ�����6� pQN7}RY_8�	�^�Z�l�h��	�
�A�@~�7Z}��m}a�#R0O��AFu��<Gܑ�7BO��+�
��?�jr� ߄4�-���p�����1�Q��.e�B��so��{E�[V\aV�> �l��6;��7�ܣ7�@��H�U'����!]��w۩�.���(�K?p��I�5�+��P�Җǚ8;��Y�vjQ�?�l�rF̟Q��`=��]���	��l�|��	jv����h�N�WLq��$��q���9~z�Q/]��.��Ң~���`�'���E�븶m�fgS\%y�Pq���XMlR���UM��m����Ɯbyd�7(}u3l�'��R4�wq�l�1����4(�"%���,��E��%F.<�.3s����ܿ&/!2<�\��$������~���)�~QN��Ȥ��F7��� ��Hu�~`��@��,1��~�yG�dgg��43�BV�M���W�y$�-iZNi)�;	hy�V�{��x�G�Gt*�_���Q��~�M��Z��T���v"n�/�à��qd8���O���/j,�n��u�̖�"��|��0�� ��T�I��࣯���r��$�jܳpZB?�.����zvJM�Wc͞
8^��Q� !-�E�mʞ��'m�Ƀ �}����{ţ�.����5���a�N�3<(v��.��qWF櫱U(Z:��+�['�,qJ��ݽ \���N�v��+@�ɜ�hq(�w�iDv@�Z%G!��q���_��ڨ�����ծ��b�A�X{b��q�+Y<�J���)�Uq��i�;���P\)��*r%v/�ؗ$Մ��{�+%�����P�W����bӔ����U�ID���&&}F�p 3 (���=��7^�����B�n����L���{?�X���t����[�+��0�ѝ,�+��}.g��;��N���"K!�;5֏�K�a����W��!������`f�RXo�O���t��M���.�5��ͽe6Y�Y(�����L�8-^qQ�|l���Z���r7�K�%��Р��5��PV�F]�A�������"����� �g_h������߷y�}XB�Jɋ���Z������3�F|�(2�V������d�r\A�=�6��W�`+Sr�ƶf��xg�R���q�|0�P���Do'
q�_-���Z�+[w0�6&��ȍz0�$�����B�I�7��H�2H��97
;��⬲��Í��Ӑ�*��/iITUr�H�@�hF��'��7mg-��A1v&GC���f�ڊ�8n�K%�d���K��ƚ,�t:�)Ѥ��A�� ���3l��0��`m��u�^/b���kٝ�*=�W�4Z�э���wCS�MILph�@�k���%/��� &��$��]r�U������o!��S��,W�ʶ�m��d�ǵ���8yL�B|\0�L."�]��~��`J�5��#!5�&�?�ɻ��AMk��A8�~'����[��D<�I#�P�1�d��K(!3y�/+�qp0���aC���Fۋ�L��2��g|�@ם#-ǖfª��v�Q܍����p�fBy�!ݶSO�N�0�Q��;e�ϲz�D
g@Li/����C��?<&�+պ�5� k��x��'RDk�8�X�c��F�l�����I�j�S�w[P�������ʒ���SS�Bo;�����ę�X����T�|��f�mM5F��;چF�w�Ĝ%T���e?�{��(���I����U{Y h���ڞ�n��aŔ�J��t��c�o��g�
�0�od��Q�䫩�@M>�SpX�|� �o9�����m����Ը�J�i���
Q�ډ֜CƂ?ٮjJ\A�N��|S���^7wp�I'c�����3�)�""9�K
~L��u\���xnj;%��dU��&wf��;�y�z;�J�y%�Y�f�`�p�hy��v�s�����p�j�Hg�ƏJ�u���'r�(~`�5��>�����C���(��C\'��%'i��dTxt��7��%�hZ#�=sʑ��\4��Õ��}u Nؘ{�KW4�y��������	D9�/YŤ�~�3�J�=����Y����d�ڙ���u�P�4ԭ!��^d�p�CTK�}L�=��(dۈ޻�+w�n�\�]�z�a*�mm��<+-����i�=V(��\��Dm~V�J6IG+�Z�Fnhj_�^�j'-T{hA>p�*���~�e}.%mA�U�>B�v/��
ԭ���FB�[N�4D�y���J������#����`@�8�s�Ĵ�,ڟ�����y���?��t0��Uc�7�ќCsA��X�p���NR�B}����p�����i�X�L�d��I�s������d���$�>pn|�e;���::�Ahs(��S�ْ�ᵒ�0��i�����21v�a[�D ׀:~�,#@&G����R���يp.=�-��������сf���ڷ#L�7n�(p���)tȹ��XE�����~�`�w�5G��&M�|ܨ����98@c���k*��/�5 "������t���T�+����ia�8H{�����!��p<1�ͫ�.b�����2[�{�+�ӑտ�[Τ�G	��F�N{���Oh���7��\�q�Kc�Ӛ�����8��Ad��y�O���A�]���q�@p�b+i����Ͷ4�Rȉf��5�ܟ���Oo��@��0���ٟFH-{Xoи��M��<��Z����o̞�s��ɋ��{�K׵!`���j�q�/r�d��XLGN-oo� �����T7Y C�YJ6�60�f�\qNf�g��T��)�mF�:M_�2KI�d}�����Icֱ�]QYcJ�J�'�Z�B���;�-�R~�'��z]�v�nj"7ب��4D��77�D���?�w���v7���)� �����mE� ]�I�Շr�j���v�@HKס^�yC�ɠ�ˉP���+����l	��u���E��{�C{>���4t%n��	"䷛��xQz.��_i�1&��YK��</�t ������|	�H��8Sg���B��ZX��\�ߒ�޶?�Qf��N�d)ǃ�H��O��o�eh��Ob2���%�x�U�M���-`$7;�8ݢY@�>-��5�:��o��b���)�L��y��Zv�H_�>}.��X�Bv��qK��[��J�徲��m�� d [G�v?��L���o��azO~�$�d���~3*��JƸ����8�( �� #�����"0��3K�rK�:�b��t�����}���Ԁ2߅͗P�fC��7-CY��`o������&��N��+�@#��=���7(��ה����ט���k��/�t�س�b������ͼ��"S�J���|^�>X�����Sq��F�#�� �Z!׮Ꚗ!�nP����槸/�_��Am��K�ɲ!1�/H�9���"A�1�y	 ���sm)\q}[�m�����£�����Q��8C!O�.#-�n@l��14�FWa+|�Qz���J�{y�>�T�&$�Ȟ�ѻV���U|�?�ɞ��c�ޢ@���%zM�|�$��	f�q���.ŶǇ7Y1��L��9��e�ݞOHo �jY Z���5���@p��z
���)�����&ae�Z�{�t��X�X�S��T���2��}�㽵���e��T�����I��-���f�)�d��x{(O���R���f�mB|r�jڞ"��j)��K�Ŏl%������Vd'5��1-%�6B��7Q-�G����9���l��o0��R���I��[#��M��c˫��K>�Kb%��=�P]�W�x�4C���r�c�`���λ�n���7�HXق�&�Ϝ��#����O�R�k�3� �2�'��:p��������A��r��őC�f�P��83N�8�րSB��`�i�T@ö(q���J�0� �b�!)��bZ2�icڌ�<����'j���猸YW"��J�^=�k�b!"O��jO�_��xbsY�p����c�	���C�5qn�=Y��k�n�t��Y�����3u*�
��Z�{�����cn�	�-%;]�ʙi[���\��c����DD� ����
B~��팒���Y�"ú��E{�OJS?XE$&v��)xP����U�#��B\�%I��bc�������<����WHS�_��=J����Z�Lü���N �'��˼�O�:@�'֢��jc� !���@�j@� .�z0P��, "g�J	:@��䌼�@��h��� RYF*�X�B��Hr�8f�����Y�j�nԁ���[dNs8��Myx������A��:�Hdu��>~n͌L����+9+3�O�T�xw�t�O17��f�cq'�a�E!�u��=�:U`����m@�@51�Ԑ*lO'�;�[](��}d�J��cj����
e�#��|� �A�_��ꢗ��F��%��)�v!9��Kܰ��U�}�8DQ�M�(G��l�gT˱��xas	�@����{u�6�7�n�#,ȣ�N�"���b��](
ue�\���A��Aw�=n*t�[R�n�}?5�������$�@�l-��Yx�=�X�Z�o�e��N�8DN4M|!��X��rO�b�s�n�52����>�laV�8�82�v�E�-Y��a�U�6�Y���v�]m�>T�����S��AqN���Q�])��A�z�q1PԲLN1ߟ�{��[ p��n������h[��t���N�oਃ>k��A�T|🱐R�gB��_����g�'��y#5�i� �LV?���gc�UKnq����Mt�uwĩQ���C$-g�~Bt���j�~>btv	�B��A�gٸ���E(��D�fZ�g+M��א�� �f�:~J6D T��~��� ;u՚����j�eA�JAᵂ���{�D��hCv�9+$7�'jow6J0;Ҏ��C2�v�k� `��	ʠ(�����~d�)�&k��N�=�|LiWlSμ3[��5-�{�Z/��>�6J�~pE�S��hi|��;LR�bVƘ>�Qģ�qC�{��W�ZJ�'�\G�؄b������Ғ؟����P�?�my���I�Bʢ�T�m��p���`@��l �� ��`��c&���='_�\��<���q~q�b��2��6Tc���8>}oڻP����Kza[����у�64>|������W�3���G��hm[�A���M�.�{�QVC�%Y^�������d�ڰ�+#�Q��
;\�E�E�s��ǿ����	�5,����q@e1BkA�j%,J:l��!�=������ZM1k����T�M��A�	kUT��@dn]��B����X��,�u�G�Kљ�h*: �=ʆkm0�0����<�P���щ�I�_.޾�2�㇙�ꈍޒ(>��G� �־Z�#bx���q�S����uKt$��<r��'4��f�#,�+z�s/�3����g¢)�Ж�.j>�o'r�$|�5�حJg*�����1T`G�L�e�@���E����sqg�=�s����r��顦��q���W��<������ $ #b���A�A�E��m8�o��1�ԍ=dD=�Y"}��oӷ����1�|bD�M_�85⤫����5V���@���h���Cb��t�0OC:�F�L(��(c1�t�N\썸v�Dc��T����O�oדa�O6�=���F�����-�N��5��t�p/[��u�p�[�z$�ԧ�6��|#t��S;�2�ҡ�"�A��}9�J0x��=��Ë\���+�Z�e�?#f?�	��/������_���A��p	/[�XQ�:D���@#��fpL*�U�ۖ,�?
����v���*R�w���I�,>���@�)�m��v�L�B�usf�
�0�>:`|Q�l��x%����&�F�K���'���D)%�\�Ѩ8a�[�9m��'q�%}�R��� cT�v/�Kj�"Hk�(�?E���BAx�Bt���1��w�վz���2��o�!���X�5-�|oL�;|.�~mEsZh����"�³E���sA6�Õ�%{]0���^R�6i�0�)�6T����n�Ets�ۖ�O޷D�D ��P�F��H.<�K40�m|��.] /���)�=�w�H��y%���A>���.h��O����^a�].��S@	e���ˋ��X[����W�tr�N&:�}GU�qc�.��r$^0
�4;�7�FC7[t����WU_��������ɲ^��q����-��k�������q�/��vI֕�@�d=~��/~�A�<+���Px�!�]a]F�9뚚�`s�j�k�͘8Pt+�g���PxYCỌ�@�^�Q�4��oT�r��k�R������/�o
j�T�]����D>1	��?���6.���DE�Sc0�>)~#Q���ʓ�h��F��#��,SM+�c�.ЁQ��46AN_<c5氚��G��46�?��q^�#�:m�G�K$6�V`~ǽG��2�/��%����ܥ�u/id�dna;&s4{ a�u����Hx�G�'��M5��|>�6UT���=u �{�ſ�Cȯ>����5f� ia������K��a,�)%V[��~�6	ٞ�^-�:ߦ������BK1`�c��t�ʬڐ;�"&�/��%ēfY�d�#�&�l.Po���&R��Y-_�2ܰ:�y~#Q� i�0[�Dxqg�z�}��ҖqY�qs�ӛ���g<z�ț����O\jL�E�/�w�����zn��W�lh�Ϳ�Zy{���<��cç$��(G�z��i�\�C�|Y�6���^VF7l�*���4UFbJO�gk���,9Ǖ>�`W����]��R6�dWh
A �����lD^�	�)��s�6�;3�ky�u�f�)��bOT��'H+G��<2��x�?}�@�q�N��k�����V���R�H�3���7Ժ�k�`lƢW^��.�Ζ��;�S��h���S��ek}�rA���*N\�|HOa���U�v���BC�w�6�!%��/�Y�������e�cO,��M���{d�1j19=��>�"Ϲ�wx�B���#s���so�1����aVa	p˲�}3�Nk��	���WF�� ���W���#�.���w�v �;HaW�]�Ar�ѡ���)�
�nyqOch���b������.�2�Кg2a����d��=r�1��^
4���6��6�2���#��v?�I�H�U�1��[-ͬ|��rz]>o/w���&��B�6�1&N`˟����P���>���:4�
3eܢo��'��xoT?�VU��������\�q����4���JYpV�e��~ҷ�|��2)��Y�᝿�QH(�S8 �!�+x�����>2d��:N$p�Do����9BU;I��@�`7!5c���>^�/WѦ���k�,0��iJ�%c�OC�c5�3N��#��C�z%� ��jh���t��_���Ő���2��~�4�H���v��B_�遀'v�f�����#�
i�iA���4D��	)�R��{N;^�ܒ���np��U���m���d"��Q�L�avE�i��Ӵ�1ɔ��=�2��=�y�f�(բ��G�ׅ�)�f����V�Ĭ���|�d�*��9�"ϥ� �s�B�0���WB�{v[��O����^
���F�⵼��|�����6�m��ʬ���^�$y�d20m���{� [�O����E��]5T��Ο#1�p�s4;��m[�Gጿ{,Cv���P���}�.X��'����j�
k���"xn��t�YT+]�%�v� ��`�K(I����q5K���o�pj�߅(@�PV2��'�p�AV�!e���[jz�Vu��l,x���Z- �NWH����!l�4
��b�Ji*����G����Cv�	����� ���}o(��8w�9����;�
�),�0"@$�ڠ&a�^A��6��%�8yn�P��ݨ�ЮN��DY��}�EhS��#���J��v^Ӕj�����~��]�m�2���Y`#�M��ٜ5i�lX�ضa�M�]f�&)4���M�Z�es_$6��?���l@ -����J��o8�]��Ey>o��P�/2r#u�]5MYAj�铬�V;��O���щF�g"T�����4���Fj�8%��tN�12=��H|�ۓKe(_�h��o�t�����Ϳ[?���|��!�����lK�AJH��c�f�wk�&�pB k~Ec��gf$JѤp��%�p��4<�I�L}�z�0�K��R�j+�u���ڴ%}��o�1>���h(&���X~:B/������6���g�;GW���o�$����OE���B0)������e�u��RWY�nz�h{L��ي����p�Ʌ����+t�;\U{z����-?�D�A�\afO��h9'8�@&�'�_����1
�-�r��I��%�veRF�suV�ԁG�j�y���`*�n��Bu�r�욜�9P�����'9X"�,ɼ�<���
RM�Y�����c�NN�Y^�5��(�.`'�Fx�
�I\!�J|�2��1W!<�Y<��H�(v���%�FKKJ�~0�k��q�/�9�7���_Er��%��m.���һ�w�jԀ�>!��콚���]|9�����k�^e7��K�kU ����8ۜ�����u���T�I2�2]�{�'���M��&��^�@���JAz��\��z�sr%/)P��TV0h�[����K�J�mZ����bM�*�!�,�����FC���Ƽkھ�V{D��J+x�%��ɯ/C�)"L��?v0������R�����$W؎�~ �~��g��O0aX��L/_nPKc��]�㉄B�BR�}T���~��I��UXB��+>��k̓��--�j�ߍ���l͟��72~�7�����p���al���l7�0y}�m�*P�r�\�2������6\**���ؠ�Dy�N��|�eC�-�]�N���Ǝ�q^��!�?�;؄��
*�ܛL2��<�&��T'�i#$g��r.#��-q �����������5�n˷W(���хHχ�)c�F��&� :8�?�*FΧʏl�fL|�Yk��	��Gz�ru:��d���]%\�8?<�5�!������擾ڏ6ͥ*H�[��5r���6�5R�ս/oeu��u)Sْ)t�
���C�'{�lIX�wA�6Mը_qp2�9���n7��c!�أ�Xp�X��q���"DyB7�H���y��2�'~��w1�/�ƭβ�5�폛z�������s�L&u8�g�kw��ߴLQnd�`�(t����"յ3��ZR[��j��Tإ�܊���
��0�|�s̡�ꇱ;g�bPg~d������>��X��"�.w�d��,�(�V���%������Fq8��1"�S��q�&��b}`G4�3`\��5�q.G���E����5���Ɍ��d�م�0e��?$��J'8��:����iav��Dm!�D5-R*�^*|M���"�y���@��M�t���l׀bf[MY�
���L0e��+���[oRF����I�;����RN*o+[�E�I$2P���4 �K��Uh����r��@�v̬X3^D"R���ۍ�y��x�� �#�:�7��6*���T�ɈC�+��5��9	;�6���nK�)��=?煝�ns4�݇V&�HK�1�,�ef�J;� �!Iz���`rҙv���j�Y1�(�Py���k��LXU�VF u/9�d#��~���.��k���t��ާl�6�왋��aA:�b��s����m�;<�b�4�ð߁��q��Z*����h�Xt"��ܑ��!sD��I/5a�u{ �y\�O?��̧N��do�5u<Ʈ�ҩձBM s�����lυ
���������	S*P���E��?�<��@ꡑ��Ei�)v��Q��De^�hf9۲H��F���?����Q�$GS�����#$@���ܒw��W۫�+�A4����/�in�4� �W�T��E���f��O+|zN1hT?�!�!v$�!���V d �S��_�yr;�[�P<w�;��Ԕ�We'O6]�J��G�I���3�́�a�i����B��Z>@߹�<W1}�ှǴTt���8�>`kZ3}�ٕl�/4\�B���{����nͷ8HąJ�Q��u�h�e��^��P�j
�XR�%[��cAJ��"_�������C9_+���]̐��HA�~]M@�;�w>$ ��	X�c|�m&$�e}{J�C�&��3ld��屆K��b����v�|��HȎ�}H���{O�@;�R���vU�n�8z 8��˧�Qr�f�`Z"y
&*��y_��s;m(h[o�{16������j�L�=[�׮�Z�k��b!�)	O.��k"���f��ֲ���灇K�%�d���/�1I,��ó��/&�R�Tb�
0ج��5 ���W&��]��U������,� �G,��_ծ���h\O��cW�W�%��i	'{M�3��3f�8|�����[p?��-EC!f<m�1��s$��<6Y��`�M���� �}�zQ)m�	��_3u�D��3�}����7�2NI��)�H^I�P�ɦ��׵B���&<�r�vAy�+�@S^���Iؿr��D�XG������c\�
�"<�j'�i��@:x\����&��|"<>��{U`�5|!_�sX{�Ȣ��kG�d�K�J�#C�]����$�y��������Fƹ��H
�R��߱�X�0�]8�Ź.�*:d������M���/�4r����z���z��ţ����68��xQB����q�����z,�����V����r>��P��m�_�<p���sT'i�N��(����~Z���ݩ?��=q��խ��ڗ���F����$j�N�*h���اe�n8��p٬}�X���}�Y��3��
!.P�
s�� 2���Բ�E��F��?ʍq]��C�:FfX5*�ᣆM:����G�N@�T�^�[�9��߲�3,�z%�����G#�����p���8[�*'a�j������,�S!����.����e�5ȃ���Вq�>(�����e��j}�ec�+DI7�l{�� [�i���gݪ���~�I�
,���c��U��i	�2s��S\�:N~UGo�{L�3#"8r������)M��&�<��HB!	�@C�9���	�\>6�qG���݆�]�c��ƫ9{S7)诠#_�#�
��D
���5���ZԠ3��M�4|T7֐�I�̜�:���ϸ-��.s6~Ę%6��*V=���P)�-BM���۴i�l�l\�~X8�-�g*Gg��Z��d����$���@��0�ܛe�J��Ʉ�v�xڮ��T��c�V�WG�0�Giٝv0v֐�N�|�h%mI_/�J��_R�8�6��
����0�_�a��"�}6��|�й��)����=�]?*�j(o�n.��H�4�j �2�tt!�����9%��m�q�>re�\o��T���!A)��*52�3�Q$Gn�4��V�<�쁩}�x�̵`h�W�}?/̜�&�$����ʨt	���S���l0��Q��h(���6���!B��&r
��f���6�Wԉ��./\L<��6� ��b��g)ո��y�[��nXUC8�KNIA'��R�B"�l#��m��*�����.�6ss�AP�^�/&��LCօ8#�ew��!]YZW�R�XAg�� ���z�'�A���L��k�Z��`�� t���P��!��{���������p6#8� �~�9)m�f�޸�IG"s^��܅Q) 	emp{�.8�7��̤�k�鶹=��hM4(��
F[9�Km�WF+Xxy�:`cS�}=���(�XL�k�*��~��C�M�6�#\��vT��o\�YV������~ 06���&��W�<|cf�V�:B����O }�f.��q_qSy����c�Z���A?+js+;��c�v�0D��N�#�B���*�4��\�Z��U��M���HǶ�|�9��m~}��'ʕb>�31#O.T-�R��r˼�0��W~��[�8��l���L��o��W|*<a��
6]^[��"�!
�)�������K���6�5��D���⭟Sa�
J���,�n�<��Wл����DHv�*4ϻ�4{�Ξ�)^$Ը}s��8�ٟp�L �b1a��!�eiq{,@ l}����3��	���E������z׳$��I��K+�0B ����L�W�f�Sq.yzۓ���/�ψ|Sn���k�ا³ǔѹ�
�`�� X�R�4v��T��%7�CT։�2�f-�Q��r2�^������GаI:(�.��Q7��Z�}r[k
-�V��u��n��\�]_X��;Z�/2x1��(EQB��'��S��	y��OF�G����mO;����$����$�|���Un�o��Q������(�V��̖��q�#Z�c� ���p�D�i�P)E�M�P�w�H�3r٣?�Xh/������yFr!L�~᝷�b
Kb3޼�٬Ԋ�������4�WH��*�jX���Du���^�F�~�9�����8D+"��+��#�T�ή�D+�"�h��t�}�+�#�� �S��Mo�"�B}*�\�[Wq�� �
Y�W"�m6@y.��=kwm�
�'Z���	���{��F�FHB�]�I��)��}�}���scZ�2X��_w�@5��@= >���:uk:��$�Ʃsc,����.���>�<�K�to�ݏ��`����jz���[g�e�]Su���CN���|�#p��gA�c�x�ͥ v?���j�1�s���dI�;��Z����9W;�d����G���-�ڵ��O�%�A��"�e>u��������K�:ء.���)�<���NR͑�M#��Ѓ^�T��~�g���Y�u"�v��Xҫ*�U�s�v)J������(�Y�잶7L9���d��să���Ғ0�=:�s5n�~3n�˿��6���Z���vz6�iJy�Ht �����������q(��u��&.�>���Cr�D&�6S��g0A=߀��N�%ܢ�ID���K~t<B��� z�ҲC�=H�rE�j�Kj�u���cfף�z��6��"�`��kO�iR�)����y��,,ʜ���K��f� �g�BNOSJBS�����x
�3˦/tA�S��x����n�tKo�:ý�ݻ���(|��~����M&}�%�O��Q�Ď��E�U�rF܂��*�elN�u�\1�-W-����N-dr�:{�%-���g���k�i���,��a�u�8/U/�N�`��n���3�Fw��7�xI�Z��[�&�Rgĺt6���K=U��v�D;ܫR���h�R��Sd�%d��x�����b�y�;��z8�'g��o ��]#�y��i�h]½M�"����wG�;8-��rM}Y���я�y+i��`��R9&�Q��m��0���wA��!��֩�xЙ�Nn�Pr��Nu�b5y���W`��D������9"���-۔u٬ܻ�v0��qdjW�V{k�.�N����g{m����ΌF	����Ԉ��($�xP�l���b�7��$}q�PӖ;&��tْ ���n��T���M����ĂF	+�F��MXJ�!DqN���]���)�Rc��)T�/{���R�r�!���Li�m�����$�q;7Zߜ�2�~���L�i��I*֡�n�N�C�sEa��H�;*��8�V�3��o+YOì$x?�Ζa�{�U����@Ie��ղ�9酕Ë#�G�*�lp���ձ6�S����}�[yY�D=�KJ�\�zrJ��bA�h0���Em�4��
�}̢h���MS�-wSM�W!=�䙿���V'��^u�{���@ �{�/a���Ű��z��G�8�d��M�ڔ�9��sAP���M!!�{�A`iX�<5s��|����S�7�,��[L�s�n=x��ƭ�4�C?��9b�G��@�7�����B]���c+Pb��}2�|� ����t\�Q�w\ln�%o���7a�f�AH��+΅��x!��OGX�"���,
؛:N�Y�B@���B?�TR��!�Ӄ,�Z��Г�$�^��B�_'XG����L��B� �����?���]��Eh:�XDAU�	4�Ѭt�2hv�.Y�'PWsN���E&��I/霏��@�n��r�FN����ih��CTIz��A�<y+𐪷��-m�S�afP��J�K�y��p�~@R�%��f�ˤfǲ]�Rgd���f��1�NV�\�bT�ޚC�������o|B~AC7�L7V��=X~|NA�-w�f��|�?�\���l�%�l��^�ܗ�j$Nx����E�8�^�9��-��?�?��Ҡ�w�R��� �H�W/���j��1��Rު�A��u���<.!%5��Y?+vIKkj5a�-�hl�LU�\��ށ�wwኁ�d"��� yB�E<;��!'��'ȉ��*KG_E�t�M�x(~��u&��d�,"��Aɂ׍�rU����?ɧ�6&����$A��B�>�NU�BO�+a�t�Jv&A���~��=~�)�����B�%��wn��ކ��&Q/A'��g8���6R�H�Τbp�?RK�9ḶZ����*w��C<}��Ub����p�A����+�L=�Q78�5��r1��-��2ZYa���s�7��8�؃�@^Թ5��ˋ�?��d��VN=��YI�����[�ؙ���(=@��mQ������2��1N8���Ä�^�X�g:jA\�� nl����M�#Ͽʦ��0�fT�S���;;�����(a_�MPP@�0��x@yt��S�Ē�������.M���*�X��)W���>'�}���S�v�e{;Š��uՊ� ee"��-��Ѻ���,D �n�a�߆Z���ٙۮ>�##��Ww���^�yIO3�����Leά��I��S�hR%�p���J���Yh�4�������e�e@2�*{v�����n��wX���$�,�G&�<�_{�y��j��Z�5]w#\�����o�Q؂�)����h��f���i��]N$c�,����Iᘣ���T����E1W�.�����Ԉ������i:�`A�ƍ_��(�Ӑ�������Bn�9�5�="���W���:Ed���ߜ�Z��	6ϲ�� Ԝ�`&\�iϔ�y��/])G,G���3^�I����G���qk�e���ŏ] qE~�Ō٦{+.��~}��^�=�{QM���[�|۟��[5��"]��C���9;l��Ii<��\&�d�܄h"{�H4ō��d�A��[�7Y1.�4����d�|!�i�Ά.{�O��@bf��o2�	�\����[K��2�%$�z��	҆/��p]�!�L���]X�}�gԨ�\	�Ҵ�Fu����c����"34��	�5��h��Q-6����a��Z����˹�:ג�G�;���R����N��)�@����c,������"��O��c"�Љ��dM�6�!	��������U줦U˪�7ǚw�6���i�� �(+���<�k��N��ݩY�V^��l؞�
�`L��N*�h����O�`;��"�PC6YLfi��3#�#�B����F1u��1���%����J>�J�[���A$����<}N5�zjBlQ֊�����ϑD��"C�.�Á*�=��G&eB'��˲�!1�T��{�u�R�Ζ̓c�&@�+R��FP��g������PP�=��b4]�mC��Ps��X�"M��p�����h��"�g��o�E���OC��Ξ)�W;Z�������p��b����� �͠\���F�FHƻybT��Z�>g�u%�����(_øo{c³�����>��rP�؀��=J�ff��Lɓ;��Ke��t���r����L%��C̒�煖jHp���_QZ��Y�-z41���S�y;芊��h�KE@r����$a5��t#Ų�Z �Ee�ς䉁���]|V�,�\!��c�!�"���O���N#*1��,6�v�#���U1+�}F5>2��7�ɹ�mǰ��˙�HV���u⟪Q��[��|ɷ��!��&��_�O@�#�4)����}5k"�/b[J&�dO����t�Q�^#���3jFK3򂥗����O��@Q�Uh!Gmu�l�����Q .����'
-$�gdC�Z�vo�~�d��v.�aI�VW��Accȏx�n@�z���Ļ��a"`)V��uq%Db��¹֌��U�E�-xkHn֌o�I�-���f�NQ?N}���>0M(��Њ�C������H6�BF�)���.�i���#�݁��b{��@�w��S@��h;)��f�{teݸNU�[`EIU=/u�/��׏WO$8��ٗj�w�~ք���fQ	�F�
!�>���oP+�J�_�W �t��1�ˠ�z��>Mt<�;6�(0�A�<1I������j#LQ����`J��\�޴�ݍdX��{���v�I|��p��p�Ǣ��3���<@`+N�T����%�)%�Rfԙx��V�����A�^MdO2!��՘Έ�I	��V�4��~�}�-]���L��u�^���Z�V6�	�ٰ�,��8?�T]'��mۣA�"F�F�4E:��?30���w��Y�y �����7�/
u���#�Lh{��폝�fd	=�+�Դ~��Q8t�g��[�+��o*7�J�%\9��O&S	� B6LR��X[&�+�I�T��m n�+qK�����`@[��
Ha�2P'�N�C�"8&�O�/v"��l9��س�V���уS�vP���.S�fnI$"���S���H2��d
�aqCD��-�Y'�ϻ���o���_��,�-�y�0��Y���;K6-}�� P���rZQ�����#�/�̼�a7�q�t��kO�J�"n��8��.W_N��§�M��J0��S�䅽������evy�k��8&SKl,t��FA�b�p!#��k�+���Ђa}qPJIИ��#m'7�t=�e. l����]� p&F�Е���%4��tun&0:�^S���%Ӝ	,��2���k'�$�NNgv�T���	㢠vaF���h�PyC��
�7@W��QC	�Dzjm��qTv/��H�	Má��LMtPq<%C��]�9N���l;n�����Q~��R޶G�~i)""�����"\|�DE�'��)AŹ��0-2���JpC/L�N�C�R�X�$��af�k~ UD��D���d�h2N��2kBE���̇�G���~�i�$�ܲ�-��F�}���f�]�/0��	B����0��.���]��ы�?G�ڼ�euF�.��/T�����o��Fe1ه(�(6����N&�{1�ΜG��ȹ�6��z����sl�s�x�R}f!x3�ޕӰ/��1T�+��:����T[ҭ-LD[ztF`���6�\�Rr���Āc7��R���ϔ V�Ka*�ϐ*�FU�U� ��t�!��,��O}�׽�_$�I{=&��C��D}J�̴J���c0��}�e�j7]ct�h��B�1�l�f��oT����p�� ��W�գ��y$P��C)	Z۽D�{��
������z/T�۱ښ�XܜmMZ|�k$\&��+��6�.�*�Y���N��g�!��Wz����i�o��c�O'��c���1eµ�Xb��#��M֟S�6�;�� ��f#�-���E��o<�]4��h���������y�?�d7�1V'ɤ2�.�U�ޘ���T�vP{�Z,�,�TЁ��b���r�J�l��cp/9t�Gsғ��9k��T�����2kPX�S��I.�ڄ��rE��@�0v���]�LS���"Y��M�y��H�P>5Re�	O�6��	�6����aEL�����^Й��T�F��O�}{X4�u����˜�h��b;��I ��mqW;�9����\�6%�|%E�x�3ţޡ�+����1Rһ5�Y�����}��@�x�֙� ��Ef��hI��o���0��0H�c�V�4]N0��$*}F"�mױ�HO���_
D��|P����Ml��'�x<<J��1�j�O�@)U's�v��d*�Y6!�]hf���B��C��d(�hRwK����ҏ��]M��1c�����G���c%C����8��4E��	����Z�|��ʢ�咤��*��5�AC�'�Ji����u�)�w��5�����尉;�&��Z��_��ƘJ�Y�7(�����d�1��pZ�C4L���cŴV�d,�[b�B�.]��u�|��:5��/2���͍�m	�5JGg*B��7)�sj���W3\q��q1r&�&Iku�0�_�+���@��t�T���r1=\~*���G�����+�t:"8�ِ}��Oǯ��"ao�4�����,�x��{%bIZ��3�9&����JM���i��������z�.��χ�����X�_�̬ d���A�Q� l��麙H����j-�4�&�թ�����Qv�5Q],���)�j9�z��k��`�C��z��Ǧ�[�8����h�YtM��b��n��Oj��}��Æ!�Ezv�'�H��茂�j�������
#���L\��fb�A�	���X!�4�^����̸�U�G~��Mvi�sx���6��=!�h��Ws��[����W��(�w����V��{R1�X{�h:���a�2���GJ��8۩�F6�u�;9:�HH�#�U���*B,����8j%�M4$��G
F��"t�n�p���Ma{x�L�u��.w[l#l{i��h}��d����&Î�[�%`6	�[p�X���mBg�^��w��	�M^��s`-�Fz���*��o�(�6 �T��^�9���j�.��t�LѠU&u�`���N tl�J8��h@��V��C�ʺ�j"V�y����Eb�=�h�W4'�W	=,Uh!��bi�٠�\��\�M()D�pm ��qv$��?LI��RV9@l���>���qtT�:�ˑ��IE��q^@�a�֭� �E�&p-+?x�`����ѶP��_�T�=`z��}={ne/�Bm�ӗD�\Qd5�Q^{N\L@�ϠJ��+�0AA��cL�L�vQG��rňtܟ�4Y?V��a��kaI�ZG�d��J�rT`Q�bqkW�đ"i�* �ȩ�3�k����MƄ�	��>�a���yF��K��JL�B�c�n��-��;()�d����N��S���_^�j�T���_�/Y2���@D$2#UUu�#���$�~K��[�*����X�LJ!�G��	S���*��#qL��ٱ�9P��H��8���M==,-�-�!�a20�IZH�1�Om���9��El��oS�5d�ySTUtd��U>^n�>���4<7xd���X��j.��d�,���3"�Q����G����^�0�����-�Q]����|J�Z�?�^~�'�H�^yq�4���) E�+��mm�8����n�����۲�4��/Q�)�g�ay�,��?����̫l9`i��J��A���r9n�~c�J�A�UZ���X17��}�����|�Gc�,�FGA`�16�D�Y{-�Nt��>��>M+���`�w(`�xI���zࠫ,&�Y8w�	k�K]P�|�i-s�{c'�r���Å��`wo��^a�tņ��O1qPT�O�b������ �f�";|<�:-��EYS��:Ȟw�q�28���/{�݂n�D=�ݴF�E���0xU��'��	�q�jn����27�h�kͭjoky	Z���L3iI�!���9[AOQ8�g�^�,�w�Y2��S�itڰ��"%�#���[je�!��ݽϧ>S0�o�M䪄<]�ݦiyaU�M,���};ȹ9�(�}���V�::�V���rn����r�1/x�$��z�5,@� ��:�]�������	j��݆-��E"b	�^�.\���B�,��&�m�FA����7��`�	��*�!� ���#���
Ţ��o�w��M��5��6���'w],#un�����. �Q1��?�^bE�+G�bOI���^��<�6�_�����F`='���HPᬼ�؃,���n�R�x��^im��$�,da¨��{#ڎD���)�p�-ī���;��0�Y���7E���I%�gyz�y5z�5֐�O�ͤ!�������ۑ�{#�3lG�G@���*���	�8�1����>D���P��O*z���Ci�wƱ��E�n�II"w{jJ�	l�8.e2�F��i���,����)���A��I"���y���l���/bTDeI�{���͈:��Ĭ�R�7���0�J2�0>�q�4��>���U�0�,og9y>�A�7*��4xCA��l�6��r�@t'���y�)���	�S��H���ac�J��6e`'�jGG}�Z�!�a�<#k>2?���<���C`�f1�/�3i	5��ˑp��r���\��w�<�>�݉["aY�%2�߶4��YI�����a#.��hv���AU�r�!�k��	o"�8�$Q�F��9��/�4c���ըl��G�(P��W4˅!�Kydy�4�9�H��=ъ��1�#�x#.��55h��K�ƪևd��ge����<�.3_6�y��S�to�[M��=A#.�'��o�8�k����z�w��<����(:r��_�/`"����g�������*���1ӊ��I�p/����0NW� ���*1&�R�i>�4-����I��?	��}�
��ܰ�HvEFn`�9C���l]6X�dkt��P����҈�Ĕ����?R�J�<#<��4|��w�[Ɛ���?zP?�q�@)x*�an�����玢@��:AV���;N'H���!w�ɡ��x
�y��$5�k@1ߌ�%�<3X�B&�9��P����_`�K���#|�"kx0�N(�4�we������Ur�K�6���`��`�d=�~ocLǕV��ֲ�����K�4�j�[p�T�HIl��ߪ��\�cD
̀r��O�F�'�
��6BJ��_����$��.�7���c�:����[p�,ڴ(�6bB�C����fy*��(�$��$��'��3����k�@��N��k"$��AJ���	�#>q�e�\2��Y�hh�2�X�۞�d�ƙ/�˜6�G˶���ٴ rםDn�A��G��-���mm��s�Q^���Rĥ�HR n��,%��Lo��1I���<.������ۈ�ٙ���t��S
f#[g�i0|����?���]�H��o���P��b��¢MP${n]�"n�Q��-���BI��J�7��Z����Ȱ��;	Нp\F��2��%�f�p����8��?��r:��Ѝ=rI�����7���Lˣ9)v���9Y���25�Dh���,��U���ٻ��fʳ�"�&h� k��V�sc���h�.^�5�^�e?$7���<�uL5� �T���Ɇ/��7�;�1lt��:G��)���z#�;�|
�9: �G+~��W�J9D�Z7��>���L���":P�
9���g�R�:��:!E�Y��)�V��&��_�^��Yt�۾�Eeǉ�C����tŽ���|U�ŲN顾�����
��_�m�6�L��l	L/�����bf&�*�ƨ������mrf'��77�g4J��ծ���(✛�C,b(R�3������(q�>]�6��	��˿�{ģ�J�f��B��J|<���1��T*%J�7�9�n�G4�c�����?�f�~L��!q����V�}�٬��t��� �e�XмmI��Y*T�C�/�y^�M_�\�Cc6�!2��W� � z<�Р��d7ݱʶ����Z���U��O2H[��H��](;�M�ʆ]W�"�)�򔻧Y���(S��x�����GWxk�l[�>���`N�7#�!O��W��V��W>�jѳE�f��P���+��~fZ<�[���[���Q:qQ�K���e�Y7\�&&%[�$S=F�L7z<G�	٢�rZg�C�a���*"� Q��te~|vU�*��@юI��W1���˥�i0�����s��4��N��,�њ�*&\��Y�o������7 �����
����2���%t�� Q�V�Z8����� V�rΚ�P)w 9y��/�����;V��~w0�y�f(��K�K��\�9��j0���������m őĻܙ���+{0d.+!ɪp��uI�Ȁh�^�p@��ܻ.�c[mB��������IYh�1��a�Se���f\��#�Ȧ���us��t���>�G,�`w}=h����+p�lO�H�I(���
��'5�&�����e�72~�i��=-���Ә8�?���2�?7H��`�3�(8��-qM��2���?G���&�	����?���&���;������%�Bc�W
<��뉹:�"fQP���$Nh�h
� � 3.�W��{|g9�?��c��+�����4�f��B���K��w��Cy~��)Ӓ�~���gO^X�k�'n��A�"�'�~���g/�8
�x�id⬓����Q�L��Zs���~nC׎�'��4�ީ��eD�1�O`W��:Ͱ�����0�%�J���5��{�����5lg��f(�퇙�%ɓ�O��*� D�rJ��f��V���U UR:}�����Ϸ51��#NK������^�����@�˫�y�9TE�m�ý0�w[y�HU*̸�C��d{.�$ş�?���ȓd/�`}l�+]�|`A��貽�$NC���飌�̫��O|�=�ҳ����_�W̤x����s���m-��K��� i�	��SE���+)��e"��2���<��7ep �2� ��3M߂������L��r�3�vb܅����Z��͛Й��W��s\�]��I�P	�۶`���s����J1�`-��(TƠ$VE�7���o���DX�>�]ŉو����$meM� E	���{�s|ܷr�Az��s͉�Q�+|��؇Z�!�3� �'�XXv�l��C<߽NQ �}�N������������1�)�H��E�:����@2T"+mX�-�D��~[�G4�Q��ʏO�~�����8OĆl�_2�@t��be��W�"�w
8[_6'�)|��3kV�����v���P���9-¢P|�;�f\#��!�c�4����o�J��"@�P����R��9ze 
Ԥ2�}���5l]!;�|k����<�;#k/_�u��hf�bd�����v�35,�z�{����d]j���DJX@W߉�%7<'m�E��-�̭��E6�N������j5�쥺B�s���(��	�MV@9r�gZ$V�7�Q�yb4w�vduT0���3H_-H�/+V	�����޲<	Kk/
:D�˛YyÒ��I��Cnd��8�{�t��J�<����~>}u��4���' F�K��**͜�N.#�F���Sp �;���I����67yAs$�>�%�L5F�D�g��F ����`-���@>gCC�P��]���x߱O�
^�H<��!�b��dT滆M&I FYv�?n�p�����х۪tF��b����}�Z�Ū%�Ǆ@央�����!P���)M�� ��	q��6�&0�h�,-���V�+@��p���<�,�Hk�}�NC�Ƹ[R;�3۹� ����"�O�z� �Ղ�X�vyÈq(�JDFS�1JFQ����qJhZ�F]���.����6��������G��W�r�D�J�S;��d\|6j}9����%|�#n��uk�w�����ym����$)ㄲ����v ���PnR-�Gd֋�s�Qvʧ��6䅡�;?��	���t������u�:\��	����H��}Y�J ���p:�ۊb�`~��b&pk��������x�9��#�oB�t�-	��.Ϻ��~�t.Ҭ�#�g0�փ
h��	ӈVh��+��r�ȗ"�^��Pz��i�(t2�!�·��0�a|D�Ĉ���qsS:���؏��,�q��0��e�8����I��9g�B�s���F=�z%e�!2"�@^����LO	����<���52g��Ͼբ΁}pG8l颚����5.���B��6�_�'�H'jY��?�(��r�f�BJ|�;��/7T1fP� ���M{����˴���Q6�P7K�^f���-5-fm����iX��l!�P�6�.j��[53��Ɨ���sǥu1���
i���')��7�'�B�u���R��M{��g"��v���nI5�E����T4|+N ck�јkȾ����1'�����5��F)A�(�(,���o��NE���U�q��1�,%�g�~��z\������a�`�_-ѵ��u2(r4��h���a�@������
��#�-y��:k��a��Po�$���?1�^3���Н��-��S�ӛ������%��=�7�dd �J�9B�YXt���N�I�v�i�\�-��iѝK��T�A��ie\�򚸷Yb�G�2�Z�e+�W�Et&Q!>��Amj�=y˞���������H�%��w�/)�L�,�;)Z���$_��96���)�qN��_��o1��ŭE�u��%cQ����.[h���#W��YN���E9& v��v� z���ޕǼ�+ȅ����:+E*0K��;���{��52he�".0����S	���r��v���d]��KT3��Ԋ��p�Jm�?,�G��JDCx?���Sd��H+g��b��;3����]�ܣA�o��C4�*�g�3o5}� ��9�����B]	F��+J��&�p[��jp0���o)p|R��<֘�NL��A����T7�� �͒;k����K��O�5O?%�L�<����&1a����^a#������
Y��fp@h�w�Dk���� ��H짤�_{(�R����w�>����
�TL�[+�e��U8�
���R��{��UCB�Â���,�М�X�GA�?��e���9?ځw�!��q�ͱ�Yl̲����j�  2c�[�J� KUʖ������_b?G��~��uͶk�6x���eN7�U#�&���'�Y͛�y��dDߚ�� 
�rK:��Ť�)go����j��9!����l8K���ײnq P��F��5�x��R�.���Y�Ҧ�
�|]�K��,�\ģ�d��0kc�!�p��O	���[�`�_vܿ��&�kl+9N�i
�ݳ8`'�:C�n�.
8�-|.��H��m�;����狡����\!b�ٸ��t�-�S�D�S*R���?z�{�g�-x�� Y�ͮ��|c�7�m=����k�C�]Q�������.���i�]1#����
�PTr��n�����{�"]�\?�x��J�&�k�Ev#�
U��G��E���j<�����1���π�������br���`3��j&7QoJ )��#��Ŕ>��5�b\��W�0�ј2Q��j�A����qFo�!8�B;��R�fd���Gx�E7�Ȼ'	������3�-�8jSۏ?�_+�G8^!��򔉁�pk�j�W�`��*%��+�<D=�?Ja�G���8g�C�w�)�*�J^9SDï�;��������އU���T;r��'!�Y��`Q�a]> �W�+�P܋��6��G2��O2�$=w�"s{���]�m?H���{��*��o�qQ��3��U�)(7�17�S(�#<��܉�U�8 �����������,�G�+�4��G���������b����)�%1��i'#��w{Íǚ�~�����£.�ih���#����n<�a W��ֽ�Ճ�m�t���
��������=g0�����e���σ�^�z���f&�O���|<3��M)�Կ�����ե������>�s����s�uR�e�����[0��_'�b8C\��״��K��0G�*��'![ײU�i�$�
(lP<#8g)�%�iw2V��T�����!
�U���*߹��p44[}���s)E�#d�o�1jۉ~!&���k��>#��uH>u�ak{(~<ۭp���d�L�4w�>g3Q�ؐK�g�3K5�Կ�Afh?H���K��Fs��	@l9)�uN}r�/�T$R��Փ7�v�d ��l+[��lb�@�ɼ�Q��@]8\)k 4�t���5`(0����ǡI���d]��]�Gȁ��𮢪Ά��b��M��H~F�D^װ0��fzk��ZQP�k���"^�Tݤ^ �+�L7R�Cv��6�͓��jW7'���w������'r�J���E��t��$�!�jN�Vڎ��f�ᾒ��o]��Z�z��i!��]�9������xno:;Lg�0塨M�I��Pk��t����IB�� Č���6h����e�p��l��/�sij	�cXSv�%y��"3/����R�M�H��k; mk˚�ts4�` ��T�EK�5� �c��^�2[�}�+`�gv)}���dѬ"W����V�>��G� ��Qg�ȭsm�=%�&ݱ�nm,���14���b��)�9�p���=U��b����~��j�-�.�>H��?�NzM�#�b�fu�2��O �)a7�ż�	k��T5����@oKR,=,ji�O�h���J���Q�z�1�-b\����}e�R���ǣ����Ψ���UQ~�
��O��݀�f�p�mFa�n䍎.�&�o7�Z����p�E�?57�:I��4����	�6c��Yv ���E��'lN>�ܲ�k�J6��}CN57 �0��.:�"d=-:!+"h�^��=�N wC���~��;1�����6�ƽ/,��OCE@�+b���A��y��!��fr�{J|��޳؆��E���<=��ً���أ��Mˎ�u%&v3�m`�4��� ���ե8�:�Ŵl�S����*|���y��P	/���ھ�H����2g�/�>�t�1*J��^�������Um�����$Dy�/��7�7����M�@���_����Ă�++v�,P�4.�ԎX��FB�������c8UJ�Ľ�9�UG���C����p���m
��Q�0<#n�D:���\{F�'D�n���kB�ez���T#���G�xL.kI�i1�4���w�v֯�Zh������PTD�7���X�y/s��
Y.�+f����Z��f����	fQzYmt�{�;|�D�F ��%��A�������e4a:kP�>D9�i�W�,>J٭�uȄqv��6��U��e�3�I:���N�%��ʏ'���Z���w��N%%.��	#�x��<|W%�҇����!~'���>�sH�@5nwNƋMM �G�^���Ml��S�5%��!G���>��j��X�t]qN�aᵞk`�i|���e�P��a-u����f9�ѧ�<��sK�#r�.F48�,|'�A6�(qfIز3�R��
!۪^�:V��6� 	��*?Q~d�J�y�X���x<�Ry�Q͡��4ir�z�s��π��k�a����6�&@SC>l����[��k�y�j�l�����*�5��<)A37�B�@0!C���H���10�}�7��Y��^>�������V[m�B�MY#�d�if���p�nq�*�q��clƘ��O3H�	�+�D +��#G¨������(U�>Q)��ο��a�]�2�g���|��r1�x�!�N+qϾI�2���!�.Fo�P���9ׂ�C �<��;Ux�V^Pd㪛��2�,՘WH}�������=A��`{�و4�d�,��{��"�1��N�Q�2%�	&�w�D�[��>�n2��4��
&��Z�&��g�{Y���[N��U��@|��ֲ1^d��6��f�@�g���g���_���2h���.��7��R��5,ehoY����Kg�(��֭��ڶ=�B�!i9I`� �п���]���h�f�{��`>����Y��i�+�c�5w�vq�:Q��y5ٝ�#*�؎�BPv��O���z#p�p��TY�9�8ʳ�z�GG?����@d�ugk�)�6�\�v��� 74.������77lov}����k�m���L<�u�ӽ�&ad&�s�1���ɏ�6� ���D�6�5��p5đ �
H����ss����r�1�3�����!���P�ؽS���ᚍa��VV���ڹx9\ ʬU@�4*���l��(;�
] bOYc�I��DO��#�[W���F�(U4|l����.��';FP��7��4V=���qQ�}��`a:u:)�7=���F� ���z.��x:|�	���Faj��9GF���fCD� eJ���j ��h����tN�2T3��j��kS��o�.�#˒��3�Ω�n��A�u$�n�n�-��C�ŗ,܊5�a߂:5�H����E����{ �����i'�%�[�/X��|��{�Q]�^�HZ=�%��߅\��;+��&���^���n�ԣ�7��dB���>�������S��R��`���"J���Y�%��)����]C#�5�P�z}	j���d0͜W��h<T�g�;T��ϥ2 L66���―P�N�RXNB�7�Rڼ��'�n=U��r�0\������Hƫ�)\�������k"�剧��J���>��*/qP��}p�gM�JR��������>���E��$���5���M�
ě���ף �Z8z����d�=�zɎ4�\4ԭrd�7E���.�:.�?3�n 1�����k��uG;Z��&a�o�˥1C�6�s0����~eZ���ɩֶ.�B|�8/C	��OQ��*%�,	w�s���h!�a⌿�2�]Ԁ�ӶQ���1���r892��ue%�YPU=��&li�i�$�Y�~[5u���?-�^��h����D����BHa-O�[6�6�w������0�"Yg�wsv3�l	A��܅�����I �� �D�%F��jN��|������
�L�<&ׁ�4���m��BeH�Zc���v/Y��۶n��VN*�h~>~u�d��с�	�I\��C���Q��������P�#��Æ���z����fR[�,�DqyE��i܃�<�_���[�zGM�p�C����L~�R];h���;7���Oq��5�R��;�S�j0́/��l������_�]˫Hc�%Ȋu4�5������v��m�X��C��Q\~�#xg� [veYwq�R͚$��beD�[[V���錠�j{���� ��;�qo������� 2���AB�4����}!�������t��aX�Y�)��3iR�x�p���=sO{���Vj�L�%Cȃ2�� ��{i�h�[,F�ս֍�!"��&;�[d��"�$�WAf�I�i��:�zLL����ڬ�Dֹk?B��NP�_�r�Θl��t�Q��$� �%�g��򗅳r!��HI�J����6�-.���K
E���+��1^�M�w2�7��`k0�8����R|I��K��f�T��;=;|ȞB͎M�������3�U�.4"Ӊ�/'~�A�ukT-��P^@X�5������8����`<]d*R���x���q���y`oN����t�&���Am����8|���F�=qkN�b��w8�V*�k����u��#!׸ڬ��"�5-#R�-}�ɏY���WW�8�8�b�����$���E��<h��c[w��֯$�!3�{��[���f�`��ʢ�n�[���4Q�wS��G3�<�HT��Х��)�pQ�
1n�x�&\Ň�˪����/�'��rF:�y������&Mӏ���䤩L��6�G��>L��9���|�*�o)�h��J�A�ԑt�^�3�$��Ȍ�O���`��py��\�xǭ��H�	n�L�D�ص��X�H������I��Ru��%^�6WW��,�i� ���*Vw���AJ�E��XC��j��Xq�]f��<Y���&]l9+�8+0�����Ѭ�>p(���84�@q��m�nT���aZ1�3E�� 1+ ��h���c�׫�?���c
f&FT�c����˞y]B�Q��Y�h�!n`+�`h҅���A6���u14����T���C�<n�F_2&��Uˡ$��0<qo���_�����wS�RI$�S�"��m?G� �����ƺ�[�Zm����kSt����� �J.������'YF�?�Jg(��i���Τ�8�[6&�!�y�b�'7 ���F��>�f��h�^t�����`c���c¸����\�%!��~U��"�URE*H�&C@����h�	1�pG�w��#:�P��0ģ��l�}fæ����=:��C�Y��0�.���6��C�zQ���ڔ��N���8�]3?�}�s΃�vk����;����ϥ{<����>�Ӡ-NG�o}��O`��?/�U�J�����<a��NϷ>NM�.�$�Կ�B�v����E
>2?�sP��Z���7�<".��ae�VD;,,���φ_�o*��y����:��e��f�A�nD����a��&=8�	jN��U��fb��*��&��ʞ�*�SIEm�ݏ�-oo� �f�9��|2�r��}X�iEn}EpI���:�<��u� C����H��OP�/rkݣ��[�{T�;M^>��cZ6�C�d},��ֲ����I&��Rq_�����S�O,p������ON:���/s��T�ے��
���!��J�C�,���%�1o��05�O����^�b"xp7�iY�����g"������~i���c��m��iP�6�^��T�TX
ʔ-o�\��R�	zΠ�Cń����2}���
�Ҟg!�U<������.�j�>���ް ��S���·U��Fg7Bg�f�X�R߇a��{�VR�a�I�P�"TZV��91��=�.�/5�kU�~:x�����-:j�Ԛ��N�r�g��iXe�]��/*|�](RscJ.�Xh��vr#k]����~�m����^iWxfq�6i�JJZ����*���ߩ�=�9@��i�A��v++fk�rɪS�x����f��l��L$����0-�v=9� Q;� {�
�O�RD�j;Y*�^ش�x7�����d��ۃ5�@��M��
.�����D�mHB�	%��_Ƈ� `�dܥ�h���s�g�P���F�����u�ůlU_u�D� �g%��p��\�0T���A~ײ˨"�bG�D�����ԍJw��;�a5�DlN�� 9�?���i��~nM�1>�O*�Ep�&�!�4Jz0��OD�a��=a�o��rd��5<I��l����f�'Aa2,��U��P���{�J����pm�hE�w�\���4vH@��tkv��/�KK7n�.Y;���Bfx�Q���;��j,]|Ѝ����z�vt�y��#��k�&Ka@�ʡ#
}�?/��	�� ©�I�[U�XX��X��H����r�x�^�v��!@TA�-����+�aȒ���@W>��Y*01��u'+�1�G�;���jA��r9K*9���)�ď�#:.�╴{B�ݮ9@�E����[��F]��>F�7�P�x�v%-� 9��烆.�n��)���2nJ�aá��ϑ��Xf��8^�^��M�i��8L|s�ׄ���=�"��@V2Mp�j	|GD.&�Z�@4��$�v����N�B��uX�~;���
�����G����q��S����w�L�H-�,����%!��,�R��h�� �}���Kͬ��?܅������H\�e7cDk��Q�0�B�q���tk����i�KX;z�p�n��\F�kŝ�ۈ�Vzlh3��]��I˅����� =BM�-&ٔ�Y�
�� GP�l��ţM�E�
���z?=�}⢽q|��f�bm����iz�]�����Tc�] �s^�6f��o�"�_�x��㏜~�[�5�&W����H�u1۵�?e��B9,� >���� ��Ȓ�H�`os2��ޯ�ɩ�KR)r��v�,�.�)�n�XO�W�0Uk�CT���ճ�]��Q]?j�I�v�A��N��ƂL���,��A%^�!wk����>S}�o��''5$�7Ќ����&��'��S<gB��S�p�.^kx8kT�
�,��Lcc�&H��r��2cv��Ǖ󍒀����b�,�FA�ڜ�T��L �#9�b^�C�� �+Q�ieCh2^��%)*M�g�����JIjB��m6��=|���3,�Ҝ���0.uu�y��h��o�p
rE��ƹ�0:kT`h���C�
$N�U��y�����In0KФ�ө9����)e-�PJ�$�l)%5�����$92�,�z����x�h�����I-�%�LbO���G��0�Q�s��i�xr�<\4-x�j�[�|f8��3bi�\��y���h�J��r�]�d�N�2sk��Ӈ�[��Y-���SN}��^t�A����Xs�AƠ�m9[pJ��ƜL�z*d�k�F��~5{²���%k���L��o?&�!�E,3�������	���pч)p~H��t\jrl�F1R�v�Ǿ��V��eL�	�����,��̄�𿦶m�+���\��E�WM��҄O��o@^u۔����!���� W���1�[�����G���}�G��"��ʈ�ǵK!��Le����o�HHT\��9>��KsV���v��%�� a��([����u���8]J7zC��
J�:�A�����?Dfӎ�'��?�,��{��\��H+�������Ac�BM"�_�����T�Vyk�: ɋ�V�ޭy����ԥ{�╬kc�Tk�٨Nl����P���5~+�ew��g:��]>����E��7�'�����c[�s�TN�j�i~�`�Ha�I0����<]|�u8�96������@�AmM�G:�@0�|5���.�[�,2^�mw{�=쑩���I������< ���oX�p�h����Z�(���!����}���M�����)l�E�ٌ0/�$���)��M��Sj��Մaʝ4@�Р�ԋ2)Lr �`�J���'
We*���e2p�l"�!)�Y�x��G�DP7�	?�[<�R����v䶏)�Y�u��`�k��Z�e���]7A�$O��2'����>*��A)�Õr�H�t���g?�`8k�$MK���	S	�`fA-�\�_8n��y���6t��J9�6bjLN���s��Q� �] �03(r�r_��'ngi�0�
���~6Z� a�ocuw��<�A��n�$"f&q��� ��?�%�5
��z�c�.��XV��Z���$�}rP�H��1A�d�pV�"yv�[�Jf�����gK�1]˔Kt�F�j�w�S� N(�Y$}�s�Sm�|�cVَ�P���8;"e�o.�K�H!��Z�;�MX',�C���v <(1�����n=s��Y���[��R�G�$a����D�D$�N�r0uf${y^ r.ZҡK�uu �5Uu9YF�{��2�Q�($+�-ؤ�����Cm�MK~},.�J�B��)����2�*fd�	��M���c96>����ft٩��kj���*͙�Bጪ�����ŨZ��[`��4�+��"8S���'
J=�M�)�G��-�iU���PkM�4Q�1,�'9ƫsSk[�M3Th)Vtx�Й��GӐT�x+�~�O�����^v=z�%���;W�5_O/��З�(�����H)np�9a�Oo�h��m50v�zT.O^��leٺ�ӦTy �Iel�r:d/�$k����3�X�*cNl�q$E�����4����OD(�q\���mk�`�B���P�8�?1���a�f�C&�*��x�e���5�n��*����+�IH�$WI��!�A�z�k(|�ދ��wU���eT��`#���'�˫/��#�_A����/�z���V:x2��W8S9� �<�s��iˋg�d�����Un�k%f�u-W�������~�k�����M�[�rHʤ��!��\����y��8��ٱ��O��ֺ���}̎�t~�v�ǧ��A��j\!����=*�Y��q0���7��*)򿊰4A�.'��Z�}����Rn��e��4��U�N���,��)]j�>&Ƭ��&e2,��4r����	��Ws�Q�4��xP�(�9`���ـ���E�!���8F�ޓ	tI�#��%�![[�X|PZFD��Z7-���aU���q6"[O�������8e�:@X�>o/��:��9�m��2N�� �� ��x��o�9z?��X���yǸ0c�*�:(_B2\���GE��Z����BG�h}6�ŷ�����Qg��
�!	�,g7C���v���Cxg}8�!���	�ӪO��[*��shߛh���d�|�1J��j9NW5���K}Z��������>�o������ŕ�H��M
4�&sCR�w��T�p��y>�:%��H��8��ri ]΁	t(�z�Bw9�DRB��:�kX�IjfM_*�%����9�����
���u[i�'��,��A04�,S	*��zb�:��r�x4�RH�C���l���>�����(ɔ���7`�O�B�y�7/�aˬ�ƞpA�	���٩
ӕ����W�U�e_4���{��*��q�
"޼�!Rs���B��臽����K'̖9w@��|��E�i�W��y�a��t�?r��H���h�lXAc��7N,v.5��h�l�lW��n
�����u�I��!��Fem�4���㱔dدK�A�gM��C�:7�c��]�!aV�+b�6R���e�a�Cڤ��̆hrj�;X��	�M�~�9��,��ƛiD��Jž����Z�L���_p�М��b�wj5T��d%+j�Ng�ˏ�Nt��ꕛ�_bh��� DQM�߀�1R��: ���N�֔{ �FC�}�)j��rZkd�`ѰV)�������('���2b���Ӕ�|iB琎�8�ђ�e��ړ����Z����\(�Ve���Tp���q��ַdQ.H\���`=��|)n���k�sw�ȩ=�\�T��G앎�P�8?U�(��p��a�}g�' r��H���("�!̸w��rk{���w�~�4[��e�p�]��M �uD�����b�_��@��K�n�9>zh��[��BS�0TF4��E�����C"��Q��/��z�� �<T{����}��Բ���0}ŋ��r.ܾd��n��}��#��c��]'_�L\�^����r��@
�Q�
�'L\��?��n��~.��C�B.t0z:��E)�#
��*m���g����DEZ�07�>��%�ys��m���ݕ�x�+٭���6Rѣ�7������X�cT����b�bN�^�/	�(x�P-^��,��pπ��*�)�4ϤX�S�����d� �0yMIC:G�k��PN}�˕}�o+ؿ0�;��
H�	h�:J�A��Ԓ&�q{�� �+�oIU|}�6�Ng�q�(AY�1S��nTc�`vq��N��Pc��ܭz�h�-,�\��^(��%��ܲ�֦��9(�����{�z��D�a�kF>���n7�R���$ubx��m.X�N�K<�?w��Tg]�.��|�ץ�7h���O�m�&�ꔒN���t+$.+��q}�%���C�Y��K�J�-[��.�bS�v�+�jٯ�Hĺ���ѷDhDS׹?!����c��eV��Ʌ/� �"�(���� ����;�e��r����Zs Y5��̌�d7���Ƞf~}��w܈ƹdYQd9�fܞ����#����ŁSg]N֍l�����q���=�kK�z��f����r�2�ή9�\F��Eu��gG__?\>�	�[pֻ�a`q�����xv)����q�m<�ͼzߩ<�42	䯮j�IV����w���(�#ZZ��yzK�`cK�^tf6҃;�:��3G��#'�8��I�b�a��B�F��X�81`�Ҝ=���l���Y����i�JҀJ>�ԭ����D����l�r��Λ�
1����F�~1�6���/�o��N[�;�3�:\O���>�[|���`�X��6���8�l05�\��.�j���o)���O�/�IS�)AНۼ�#���2�����ҽnxR'��!�#9��m��uH�q��i��B �nA�Í�ۈ!,5�����)R�Y�]�u����菩���U�T�}���3�	D�b���<��L���Р0��P2��蟊Ҏ���3�x�R�VC�8�&�{��;���/ �0
@�+!����wVg��DQ�m�F\K�hS���ژ����,��~��W�qŁ��ݶz��f�����M]�'0�84o��p1���ao��Z�^��S�<�ۋsZTոqBخuj��+��sXWc��C+]��I�ʴ�v�3�3�'���x�! l�䦖t�s`���Qwa<>c�L�	|W]�������k���Y�a�M�����
�.�B*�l�6�`�?.:zN�P�^���������$<��W�M�]~K2p�_����b8;��7�2�G�*zw=H/�=+��j��qX"�1"Z}����I��J��Рy�p� &�����,���1x���?q|%L���#N�@�b�c%C�IUOj��5V��(�8��(�l��s�q���<���H���*s�O�<�^�8ʄ)r�xϕ+�n)D�&.��8�~�!;cS��f��J}c��R���U�)��(K�e�ő�~]����5!��q�~$��M���?�rU����\�οK�x�f� �C�3����@�xBڟh�'|��-2"�SC�ޱ��iOR�H�
��>Ɖd��QHˋ��4�
S`���p�@��/I~T�\ߺ�Pj�e�3ڹ
�X���a�ʂ�Ưz �lhh��B�9�~! �A��g�
���P���؂��:�b��9�"o��^���� ������
Y�������J���V�E`œc,@t�]f��y�覣@�U�/*W�\-��d
������`�����t�>c�����#�F�I}(����j]����JϞx"��v���]vXRT�������� �_����wh��z�̼����5��2IzusAY~��Fd�Z�����L=��H��uiE�����Cy���������F�FS�F��M�هEꞝ�~�7=�GH5h'g�p�"�km��h�^k0�����tQ�]�����v
�$�K8�ß��򑟤)�4	9#�Å���� }mN����A����$�����jQ��Й1=_}�\Z
j����8"��������=���kB<���]=��pFEj���\u� E��}G8���Ā4�����(]�'�zɑ)�:��X>r/��2_D;�>X�0��EJ�S9�¥��{���bD�KW���2B;b�W&W�b�8�4�mXd,��+����O-�C��Z��E��?�fl y3)���x�,FѷVD�	�*�A^w��9̚�ϜR)�]�C�|y�4�	S���y���X���o{pdFe'���b�O�Y�`<��8�NJ��"Z��V�
8�G�
�Y�E$���,By&w&28d���������`z�
�M�D6�?Ű�C��Q�w�d ]P�H��6��ߑ|���C�"����RR�c�E�����qm�s�G8�V�,>֭O]|C�v�0�*���hk�e��(��s!�	�1����]t6��T�E��(v�	%��$x=�i$�'��!�,�����;CQ��,���ą��|e
�AQ��;	�r\Q:��mHzy�K.Ħa5 �7����(id��ӁC$i�1���B>Q����K؜v�l��8V#���-bxf[�j�m�]ʎ�tԻ��Jf���Kľ�^�Բ�5�8S���͞y+Gj.F�2<ߛ�4_��8y�l�r{�kW�������^](��n��ff|ͅ�r�Qy>���C��h��?����Ү�p�W0\�!C�`  �frH�L�jZ 	I��eE��z[_��P�ÐZr������L:a����y�[��
�w����a�	tF�7�6�ɡ��s-��h�Q"�!�l��Fh�8�LOrd��N|I%��Z�"+H	TqS�:S�%w3�P"$xMH�ow�~$!�L(��H��'}F
���1�G���r�G�*��;�ڐ��9�w����z�tE8~]#a*��( �(}+B�Lt��Lk��-;�uP-�Rrȡ�OU�s�%9���7�Xv ��G��h���z��tJ+2Ń����oyk	s�`Y�u���!�*�y �-�Lȏz��H�,3M�&^��o�B�'w�����x��%�楣��r7�����ëv�_�V�Ѩ���[���������U��)㮿o��%Ŭvڌ���fm��Vd����c�VY�	�Z�(�+��ٯQB������h&6���(�_�_�i��y�w�.�v8�ܲ��&G���zBzZ���e�������ӊFY䔲`{"�O[Q�L�x��b+��E��m��Gh�
x��w�F�:$_y�j�-W��5(��2��ҳ�<I�:���V
�p+g��s��˾�t�лiޝM�!��n�K�����㣭k%���gE&��$q	l��,Է�hQ2�
�&a 8:�~���JŢ�����IѧުD�*�xC�&��.�%��e3�<'�_l�P�.s��8��Or�p;��G�k��7ۙ��bz8�n�r��1:����A.�����3�4^��x�,�hMd�7����br��?\�l]^�G<Ocsp4���
G���j��۩�h(Җ��.�Y���Tv����f�l�0�I�5�Y���,��}��$]l���=�*��.N�Ff���&GI���5���|��-T�_X�4�C�y�h��gH�=K���'C1��{f��DC��:�Fv�IOw�O���>�D4��RjwsS4��s�&��A�R�4Ur�/�����N�A[�(z��(�^0nB`e �b :�\�7�ˇ�'B5@ن$n���tK��h΂$��"l��VV���?�b��������ч�P�&Z�t�eѧ�Qji��KRx8���䘱��o�h������٘Y��z���T��<e�㊏�
�VO/h�o��H_����x���
���{�
��%���H $��[B�g;��{U��.@&I�=ߑ8�L�D����n';{��p�=�[T����5(�q�5J<b6����>�����/n�Otq!2@:�K�vB����}�/��C���_�����L%q����W�}�|N������lx�%���R2�� .��/�;-��Lu=g�iXM��M&�z���F�[���)�յI7B�� dc��Nl;��m^���E�ft���-;�&n#��;�q�@y&��|'4M׸�;�#y�����}������ L�G�*x������&����o���S�h�,�q��֎bbaa�SJ�?`ڍ��Q��t�;%�ˊ��"-�ffp�
��%���@�ųyiӇ���i����^�,�b���6���,{�vf��j{r��E�o�P�'�~�{�r/�Օ�F����?��6nkl�!#���܂g��]���O�֡�t�=��	̚HU����W=����x/�Sԉqc7DձԜ�z�p��L>�2����X��#�b�A��(}����*��;.m�Y�Է���*ώ.&�.w�J�V���?B�X���\o�N���(,�����#��k%puz3����'T,"����{��P�{mA�*_Z�����C�N�>�ۼ�yzc��Rv�lR�f�������b�G��42z�2۔��r���l��������.@wa����e��S^��*���G��~i>�j��/���	�� DܶN�k6Ϻ�Eޡ�R�3�`=m���mQjl�Orw�}hƓ[R�FdD�y+��p�#�
�c-�v�ZU���e��j�5��He܄�Hp���N�C*Ѽ@�Q���w4�Gj�cjީ�L�c�� �Ǫ�T��?&�&i��Ё��͙� W�-���#Cn,���@ �x��z����Z6CC��©����?N�1:f+��t3�#��'(1�̑��d0c�Fd��pͤȟOT�ph�HC*;����"�$&��
��m_���J�;������q�yg�А����$T�����a,��nI����h��;���(Vp0Z5ۡ��X}��7EvJL{����x��ci�[��O��
�K���?p�T����s�~���)70CHd�yȄ����t7#���F���fD��t�.�L�\���,g�r\l]h�N3�r�42I]���G ��O�="ښd�F.��Wz�����K��S��w諡9
��?P�|�ed��t�T�ԉƸ�o�A'cW?�J�>� M�R��vD������l�? M�74A\UGR�\�T�T�P�E��x7`�cz:N�^S&Od��bP>��8.�s�XGn��R�#k�}�]M���F��a+�����_m�}Np��X�ӝ�l�~�]!���J��S	ý3{��f<�|��*7��x���	�3~()�[X~��/�&��h����%�q�?#%���j/��v}!�%�8N�@��"*��{�F�I��B$��;�CN�d<��d-r�S{��9l/+،x"����H��B){:�m��P�/A���A�hu�N�q��|��uL��g�AP���O��:뀦�cn���򜺿[Wp
�~���G�RQ���cP�u��2�M�w͵�s)m��xB<'�o�� g�ƓO�=�mʋ�J7$X��<0m������.�~ˢ]W�N^�&�T�'Q��ߕ�5�<o'���Y�N-���2��D
�Ś�>Sr�X�*�M@�r�j\\�G��*֭����`3Iࣨ9 �G#ug41��Mmc�U{�6wؽz�
B�MPFZ_T ���Z%ϙv3�m���|�*A%9���Qڤ������|�X�v��V�re�I`;Cc�6��� ��Y��Jh93����G���l�?3	����`�N+U?Ѿ���0�.e��O@HJItQ��b��� N��c���NP ����宮?�c�z�b���M��v����#���r�H�.SC1�Ս�$�.谯�����7]:=�M|����M���$V7��<w�Rܒԃ2�ɖM��5C� xV	
#��T�=��*�O���\�Ggέ�*���;X׎�c�-Q�-��D]�l��,~Zo���3���g�6�$���T5�M8,e���lh�[Z%[i�6Y2:@_��Ue���o?<����o��� �f���^��W����*R�H�
#�{��}ihj~�(� �0����s��D�!�͹
��z�~>x��O�u)�d#�QQde�t_�TT����O-��D����;�6JG��CE�b$���e��?��������xv&�F =eA�o�wLlEM�j'&�h��X;T, x>����+ܞw�iY�/��KQ8�mcɯ����f�+�� �?�dم�Rr����iV�f���V�3�x�s�� =J�|���V��.0d՚B��	�uQx����#WG%��	�Ϭ�9.zD�2,S�:`	����v�;�=��*��!+&�
e�,�&�2-&�ƪ]fj퇃Z� �2c���;�M鑼� �p�5P;r���^�D������X��A��R���5%' {{)�ge�GhN\�a��X�NY�A�#��8~�=�y��8����zgI�$������<r��E/	���%��_��Qp٭����,ڣ�r����0���e����Ґ�
�= r�C�z�:��{�D8H�ݿoA���M��R�eXx�@7M\�5}�ۤ�ݷt��������|������<Q�&�lz����i�1�(J����
�KX��=���G_����x����c����i�؅�nȵ�?}��`���Ѕ���
>l>��5#GZ���B�������φ��J'?���W���i���w��i���"�[*K~��:��Ԣ�ke�>se�o["�&����
�[�]�J�y�'��ܨDW7�XÁ��qzn�l C�S�U�M(�ϗ
 3+$
<������$��|����t�y�F�c���/��1݈�s�i�L$k�bQנ��Ӭl U�;��$M T�(䈥�q(�V�)�o�a_7�:vO��.*�k��ޏnvP"�ź�� }�e�.�pn��掚��l>���px`��cZ��"5@.i�d���R H��Ê�t}vc���qT�kmw�ҰMp�\�bɹ"�C��#e	�{`�w���T� �����_�,"7Ъw$2����� 2|HA���C�n-h����Se�QT��_Ke�Y�w�,��6L�Cn�-���_�+H�H��'�~e1�-׍�R�a�Ϭ^z��w&�
�A.����#Pm���Y&P�P#�5�����0�Ӟ ����c�lcdt/R���??�ދ���zD���_�"���řۚ�����r3��'��*�K���U��Z���8<,i*$�⌗?F���_]\��7�� %)�b5~�9��Y���%Q0?��G5x��S��!o��>/��4#F��.̇�AV�t�|U�^JN$�4=. ����\�:N��Q�9�l_��*����8ݡ���̆23�:|c���3����m��2��K*q�Am&�9}�Z\�FV�}3���}��(�ZVQ�����tƗ����>j���S]$?~|U�ܑ\�����+w�T�2c���;:"_�X��9���1��M̘#07%�ѶD�����+�~�<��]ҙ�ϔcV+h��^|3����$'<�R��{�+ ��
����Z���RH��@CPT�T�~6�!�x���~��;��
�0�S�����m�k��a�a�� )˲=�&]�K�q׃o�Hf�34����x�Ԧ���l)�R�",�h�H�߆m�s��������xt�����<e�RAg�=���0�y�'%YQ�̯ a堧	?��X�4��T'�I� ?(�\�=�9:̫NV��2��,��~��͞�T��)<����SU��r �x'{��Kc�!9���ΰYv������4d���#V,dъ��[ǗCY%�~m�^:E�C��.��C���ǚ�9+��̓a��q7��h2Tp�z�ƹʄ�������F	sqW�;���r�a�¡��nE�6`�JfL��C'���47Q�7>����pI@��Q+7��v�gҧ+D���&#��h< ����SW�(&�5�qO��[�n)#2��5��w������N'#>���q��@#�&������1���ϡ�ܓyV�ɋ���=�7G{1�7.`�7['��ٚ�`�H�8ً���/�d�Z���~�E�D������aH��|�������:��� S�x{�r8mK;�|��u��ը�ZXeũ�b9�F�ӛ��0��l$�~$�\���m�u��_=���jx���2��=��K��g
�'Q^�a� �
�[e��c�y��I{��_V�� ��I�}|��c�7-�Z�'@z@�Ii���E-C�d�0�}8�l�H���]EI07�> �U������I��� �_A̖ov�ܸĞ�a�Q���w�ԕ�稆}m)�ph>�@�������5%"��:HC��r�~�v����Q:�3�lv��lv�c=��9c4��7� ��}��t�(�C���O�bzam&��!�&˙6�A5���z��S���Q<O�ݎ�Tg��?q~���&�_�U�]�3�&0^�z%)�B\�������6�y��7�x˶��V�<e���<�-�����=�R ]s�������;4(��Q�&b>�|�↾�+���M��5��N��z[�F�#&h�'S�����@�Q�Sʮ�b����>%���d�z�Ih�f �*�J��РS$�X�X����ȦŎ�|��q�����9'���L�����%Zh�@͟�̭ޔ�rd�L���Y;���e��urMF�ۢ��$���L$$?x���w�?�U{�~�HM��mC�D�P���9*ά�b�h0�����I���<��k[v�eS@5h�Xfo��sI�Ŵ�C+����/S+�'�uS�s~R&�t�b�[�.�U�J��'�T�\�K��LI�74�Uo�%�7Z(�I#Oc��n��PV`Z�x�M`��R5�W�8�q�+Dp��T�7i�E�_���ԓʻ��#r)�����iߛ�4���CF�����?s0�o�PX�{�pg��Ф�	�2��8%�$n��
�i-�!СbH}X����%��(b��AL�1�!�q���U;�n=�V�P�<��z�휳\�ҙK��|�0;m�Ҹ�VB�ƃBl�+J�i:A���9�T>w�]�C�O�w+�j/��;��"e@0��^��P��o���H����\=�g���okI%qp�'�G�_�� P�hH����|�JiM/�^3��R�������$ѭ{�����,��U�-�,G�^�|r�Xe	,�~��^�6���3����"p+�L�f�>D��J	H�h�C�ت�)`�:��wΆ�J�b�F-
O_��U)v������M��²ҡ�@��~�4����D�im�[#Y��}�U)�m�h�|�.��VZ|���
�?��-����
���o,�S�J�um�P�OVZD�<+���0%b)R�s;~�H'�ل1�������y�[K��,�`4K����y��wlˤ1{x���a��B��r9f�@8�
����E�;�A�S({z���y _�,����9�{)���
�PN�ܯ�Dg���9?�<��ug��Je%�Cia~�x��T�sۣ�<���S�cQh��X����X�����K��^w���i+W�c� Y��Jn_�I�|�`a�j����îySf�|[��KE[۴��U��DtDJN\+N��$��NR/m��ā3�g'1f�#�\��J8���t�n�oIހG�����sI�Hx.�A}:�����k�'Wى%�M�e�ϻX��J���^�%��ٮ-�8�1٬Ǯ<Ĉ�YM����J�M8�*��)�ҹ�z-($�K�$k�"�C'�m�'Ѱ
����4�.^T&�	*Q5,l�C7@ߞ�k���"�^=�q��.<��t�Ɗ{s���@��?���C�oi=�wѿ����T����(�k���yc_���-7N�N�K�pB.|>��.��~�6�l�j�NBĿ3�%�_�:��&˅`y�#��@(v[�3�¥�jRF'<��N�!T᳾$�>K��2��]l�R��v�U�W�����;�ה�s�G�M۽�ttI	�U��M|Ͱ�5E
���E�� F��a�/�o�Ma�z��Y&�L��ӛ��vqBZk)�C���Q4��wע�=�����
>^w�+��8/t{�c6&
���G&�kbq�=·��G�~����ڳ}>!�6j���������.|�R�u���M&'�<z\�1�w��7,�G�7<Q��i�U�_�ީ���*d��}h�L�cnqAZ@2P�����Ĥj�#-pDWu��#��oS������zmI���	�A��=�%�Ə#��ǜ�0����X&4\�b��L��y���/��M%��w)�9,_�� �zh6�= ��N���(���S�D����E0EuݢGd*0�����TA89t��HG̆	K��F��QE�����3�2E|�9l��[g���.��{�U�S�Y�hF���)'��6�^��mj(���"�[�+P ͥ�OJ�������߄��-Wd��"ޛ�"Wr�'��\�Gݤpb�<:���'-�������W��5ӈ�~�� r�����hg\m�|E�·�+wD*�>�[4�l�par�a
�I�А[��ڢ7�MÇqF�cF��%��y/-���zpR?�fvF
NsR�����Q��|5����P^��*u�4�M� �(��{�蘽5�C,�>�e�0��y�:�<��	�ѵ�0te��l7N��?�ݷl!�S&}5�r( 1�J� ��)���t�U᠆�v�R����¬V?s5�.W��T�����RYe�ة��x���A�G	 s�]�i"���zⴃ�9�x���>�|�l���U��� ����_��oⰚ��5������@�N��Q�o'���\��C0��g� ��A��C�h�����>r�ŵ����{Bg�8m�8$�X^lҍ]��HK�� ��Եz|��@/*!,�'���k����ӀȘ�<M��[>&�  V'���%8m�|:�Bz���l��C���c��S�A���Ï�>Tw���v�x��!������D}�os�;H��,��M��CMAC�xoW*�W�{N4i��0�ٕ%�q������A0��Z ��CV9��M}kU���t�t?�CŨ�Ϛ+��.�n>P�Tg��������h(����� z0c?(֒<��FΒ��QыI���"�	�'_ڌ�h�2#޲v���[���ƭs�J�Otu��t���XZ5 �m�,�gn�H��r��\@Ґmi��	]�K���TD��sL߆��L@�߄�[zil	�tv�E��[J��F�ۦ�>MU�{1\�;QRU6�B��Fc���)3-#3BUFq���'?�B҇2�Z�L\
6N�Iʧ��@�d�X.:F�G���2���)OD�����vnm������~T��3��;����������f�T��c���5�{�e.{�aq?����;���Z;ܢFhZ��>�MvB�k��]�wB�]�eBФ���с�Z�Y�):�L�`�OJ�n[��;dY�� ��m�eMmWϻ|l|l�EI�}P��c*T���ҳh�-[���Y�uن�5_�������>�֞y��#w<%;3���LCc^���$n%��:�<6(`J팚w�E3C�v�l}����V*�"G�������T�%�����aKH+�jX���P�?��bK������k,���ړ�C�<ո�[!�Hh�-[����7jW���F���J �j��뜟sVlH�0ʳ�].��}�
x���t����y"��x�x��Ѯk�ת�6}:�ce���+���ט1�U+{5敶H�ܐ�,��̰أ��r	$��T�N4b�-KR��Qn7Tsx?��2����.�Lr�ZaIr�z���;i�u�q	��>+A�,��0���!\��Y~���)9
�AN/eJ}Ӕ�M�#B1Y/��FLo�a���Fw�q��b&��mM�3�Wl�H��6j8gz��#��b��֒o����"�TR��9�n�w����#d�+���f�c�7����j4�P����w��T�:�i�x�$��m�,��>7��w(��V��|\�+�/9N�O�����t@|3�'�cJq����Ɵ`�C�	-����p���*y7������ی�Z�/�6��3�ڙ��;(�hh"�j���|uV��
�c�ܸ]�L�'�56�F�Uź�yāՌGu$j�ȳ���Fb����E��W��*vgN�^��y�,5��9��I�"�����e���A��𠕉�ጢ�)����S;��0���H򚪛�o�<G��K�ܬ��Q�$�� ���n���
��&J��DB�x5�Ņ����7�IY�du,��V�XC#�y�+Ҡ�N�J�0ZY��[5��8M����Ӥ��f��o�yb=�J���SLa�{`K�q��ox��R���!��L��"%�?h<B�<w���Z���T5����o�I#��߮����_ ��p!*�Q������� ����_ۄC��sj�
��([�1�N�l�3	o�ӶX��%>�z���j|CG���nA�T�m�$G<D^l�):����	��f���B�^~�<*�S�K�b�V��t���8嶪e���a?V�&�->�-�d��)�z�df�$��,s/� �2Xe�xe��lN�K毯�������{��w����s])���/2ǧ˲�ߚ ���s�q�f�'Io�bvD�y�&'=�B�K�E\�\��T�o�u�)��wS&����x�(��d�c����K&S��]�t�1�43��Z�R�F�
�I�K�F�bZx��Q,��:{�CYX�j?�/��#a }ғO)HoE���0$!g?�ؽ�.;ɼ$?��}J��p02x-׎�e@��nSՎ��b�,�� �r�+]��o9q^Uy	@���
CE6�)��.z����'����&n8�HD�>�?�|��Ɣ�ە��c]��X���/s@�ּ�z;�M
�	һ%\�Uuό9᎖f�I�3z�Gp�
��r��G�>h�pȷ���z^�'���_���td�a�~T1�W��@���j��Q]jT�1e�2�!e��$�e�lw��s��?/Ĺd�s�ְ
�3M@`w�MJ�Q�[����w�<JX-�9���Z� ��f*�q��]3j֝�ĺ����w�pH�W�{�SP�eS�kqK�Q��j���Tb��kԊS�q�ȁ�ϰt�y���Y櫀(k~�jo�]h�h]?�榠�?������>���\�+�ݏ��8�K��{��ƃǞxk�qx7sΘ0�M��:�"n���<O~e����n�WJ��`t
CRJ$�k(��Ȍ������m0�3p{F��E~a��-6W�2�����i)��xw�o����>t�>��
�C�6F�q�_*��'r��>�,Q+��z�Z)��ו�� ?��N򾊙���v7�
��3}�p��,�g��������d�,u?$jq��pn�ax�n�[�a��,���9�|��S���T&�S���Kʹ9�Vg��>o��dpx�8�T�b�Dw?�����Ϭf��`�a�Q�0q0r�֭u���2�0;�z��OՉ���`~��Upm}\^�f�p�[1���c��G�կP���<��iy��j�~�x��B�<��&2j�&��pc�����L���*u��e�����a�)�"9�+�^Y���pAՑ݀"N��ƅ�A���@L�_2N���/>���1��,���?}?����=/�4(F���O����$�~G㝪�Zvfr̶P��T��j5��'����+y�{knT!u���͵�4��ڶ��=���~��t���IP�LW.*�u;܆6D*.r��V�����ѓ��,
��wH�J;k�RX~R�����|2�˛=�9��8����[����|ӘߢkG�X�v��y�/ڔº�j�Z0����l1͜��G��ؗ��<����(���¬���Rv�̽��Oz	����<�C�y�"1���+�R�B���L7A��Y���Rbf)�������,�X>!�2t]<����7�}�o�;�M����1����(d��{I� .*�@�ߓ�},M�~�N0󶒪�?��.��_b�����|g{6Y��nl-��*����r��4]�-�͝�Iء�=�a{^��[-2'~b�-)�E��+�'�P/;��>�%��^Fϒ�r.[�b�NVv{���w���M��vQ���B�Q�N� �}:��t�Ѯ"78y��=�D8�/��"�7Gy/�G�<�UA^,�pb ��K�a����=��*�sL���#����� Y��jӔ�*�G�ۑnz8X�\��s�J��W�-������2a^<�#�o5=���X3�=$���9!d9�9�9o��9���۱gάQ	�M����v�NQa�RF��L-�l����Ί��1J)�6�v��W�V�7[G�r:��7����5ˁ�h&&$�Q'�g�~�S6y���Z�&3�޶&�uS����x;#s�*��.�A�<��
���zּ.6,d�]j� �ݙ`r&��w.H\�TX��^��5�>0 6P-_�\:��އ]e"�Ǭ�l�B���(��0�
H0)�F
7��a���g�]u���L�m�&���:&�P�1}&��2��	��B�BH����X�qf��Ƨ��ݞ����s5����@N�6Ձ��A�;0'��~�lPe�5�<�0��VK��JVDS��*me��A�x��"�(X2�9a�l�eF�z��(h�1��U6p:���;��]U���0N�$~����zF( [GN��}8���V�T�2jei�M�Rg����Wa���XaX"Vzd���B{�'0�s��*��KJ�a�����b�������:�*����G�;�$����(���! �vmm �o�#�Z���'�DŎ��(�1�Z���%S��(^<��dKK9�n|u��{��k��Q�[R�m�V�*���>!���cիBΙ!��r�F�P2s[�����`�F�������i鐓���*	�cB1?$���aK=wa�M^�o̯gۉ<_�%]��UD6�~�o�n���;�u/���%�{��ڌ�R���Ry�/�j-툗����_/�iZ�B0F���\?��V?���R�A�)�Q���S~ҋ���H��GC2�P�H"yҌ!�8���~�ݷ�	�(j��葤�r�Vh;�9�s1f�O�\�3�0E�P%$G�-�y -M''��6����X��ղh���A�eˆ2�i-C�
@����R��}����Sr���(��wYг���B�!�K!�:3���C�%�:F�=�iq�[�c�؄eG�4l!d���+���Bj�OW�M��Q���}������tH)�Q�m����MB�
�=i"���� &��2��/��-N�g�������� �E�l���J�󹽹Z����l��2��ͅ��1c�/g�k9�9K��%۰H��Č^�-Tۀ*v�\$Yk�iMRx��5�BQ��ǐ����A�����P�{qz���T9=�ƣ'���'j?ފME�^�oT�1n�J�Tx�CM��,<�5��S��7��ҬX���Ɇ�^���F�j����h�vO��o/8���L��,��s力���ۚ�;�xEiaH|�����;����bѯI fv�����5'�t�.9��'6iq�*�Z�"��X|PLʹ솬��wh���Жhb�L�т�ȫ�QM�'{;ϡE��T��������Ӣ�6b�a�鹠@%��n:���%.�#��������W���e�x�0��������P�K����^��+t��(�p�:-)���_F/��>v?]). ��$NlPH ����_��܏DQxQ<�W�.AF�Ց�������;:��ڧ#�����?t�2GN��Ncr�9�?���/���j̩�*��fr�~"�:bs]f�.��v6r=:L��2|T��vq�H!'��<�n��G`���}!ػ��$�<��2���������k�B.��g���ۤ�����d��l^Ʃ���7����.2�X�}9jF�D)�t���z�
Lc�<��'?i��O�o_��a��q�'$ ��|d��}e巵��
��MY��_]U'��\���v����砻���k �m��B������◇�y��`��rg�ҿ�Gv��ղ��������J�Q���v���O�"-���ZY� /q�R�����H��
㧁\d���0����K[b��)b'��Zo�A����FcEh��},���Fa������ ��UFY�v����p�
��|*�^�<�����.HAs� Ϻ3۾<צ�����(9�@��'V���
B�ě'�gv�jy��/,B�~�B�Mt���d�P�t��j�^*W��aAR��T��55��r�5:+s�ʁ�Lq��z�ݾ6���|��f�\gY�#��e�ä������+�+g�DRd�;;��l���[����x�[�����\���l��������gLRiy('(��A{{�
ü�pQ�o�6�&e]<n*l�FLzش�y;+=�E@�m��8;1^,8�9����^<�i^���0S�
L=Dm�
@����@ܜ��Ha\�٣�V�F۴~i�.?в�2�`Iݣ�~���N��n�K=e�fb�8_���N'O�%�{\8��y�J�0ݔ����T�at�(.�N~*�A$9S�6a�Paԭ�?ߜBH���O����Ʌ[��Y�n��T�`������Ԑ?LN��SQՕ;��O�>�
�.�M�#`�x�y��]��9}ML Mm͚b�ʌ��ą��G�d�-s�Hn�����i�oW`�l~��i#�Y�
�Ur��`VT~"/��{�����=��<�'���������_��GY��M�W�c�
�o%��(_*g�Feb3:�?�Oklo������.���S�h�
f�3���RX[]ס�M���.z\�x�E���|�6)8!��5.��}y���vŃ��`Sz�s��(A�6n "K��K٣���@!�=��`u��lj�v�"L�R������Ae�KK$� �Vc�) VŜC�zq�!u"'i@γ�������I;���G /�B&�����6c���+��u�M��Mӓ:X�CM\
*sp�0��b?��c8pywr΍m�����?5�WR�>=($� %��]�` -- C� hY��%�-�i��Fi���[vF'b��������і�;�(��r���ڣ.���5�x�p<DV�mT
10����fTiX�o���駎)y�[-����$q�n�����)���]�TA�͙�;ιi
�%(�7�u�튼f��N2�ֵ����^��jW��{ޅXϧ��V��F��9W�f?�E#���]A�O��;�K����]�ػ�5��U�ϥ���7�8�42�Ԥ�ؚ�e5�w)1d�T� �v�d(<e���L+A�~둖g��TJ�m�F��p���`;�3�4����ϊ,}��Z{C�x3�sXJe�A?^P.X٢h���k�tj�|��H����w����ℤ�f=};	5Nm�e�%�~:��\��ۮoE�-Ŧo}����~M~��N8!���e��by���Ws��RDߙ5ڲ���I�Ƽe1l(��Ahյ_���d�,�����GY@]�WH��Mu����XGv-k^=Lq�5� I� �u��m��:�[~j��GF
"	�L������������Ѣ�`��9n ��˒����M3�Tw���[]W�5*�A �aX�,�k�,����x�R]�ߎ)��ޖ`F�8&�;	�����G"H�j򼓲A�����J �S�E�s���&w��P��2ή�qat�C������/b��i=ǫ���^��7`�Q�(D�5�K;8w1�v0���K��
�G�$����gܚ�v%4oG�[��yE����~����4~5����t7�z��|6����#�p�kl<�`2��e+vq�l�V<��3}G�H~;�؋c�Vb �n������()]È��CM3|<\
(GK�z�֒<�a;��������-Zۭ��c�1L.Q�󍢃�n_���G��F]�:Cd�����b��5�����
��~���z&Z�J(�W����̐ь,�ő��-����yƹ�i����r 3B׶1�?��?�[�����-y
�b: Q%g!��l��c6�v~����=I������;ӐK�����Я"�i61��j?C+%w/�B�#�����[-=��?����t���	r�]��Yi�o� ��J�~�vI�8���c{]S���ugEu��f�E.>�E����ԀZf�,�W�5�1�����P�s'V�y��ű�F��[���e�ͭ�9Ӡ���y3���>��7Z�9ӯ�J2[�����FtR>�®la��!g/ݼb2�4b�b���/ڠ`t�P�#)R>�v&�k�����͋�R0L�-����ׄ0=�����x�d�/�F2څ�PO���n� 8�@n�%d��%��[�	�ڐ=nל�/�Z����T�ą�K8�_�e��H�e�Y=��e�6�e�
z�i���j��#�/�����J�j�ܘF�冭:���A�)�t����rO���7z}K*�3�6�_�K|F�����3焂��D9�6.S�,+��7��<[����@'aD5���+�Y���|�EK��ں���]p��ڟ{���jX�O?������V�@����e�>L��@&P h�uC�H�%��6S�&t�4s���V�g����V#��')�A(�R'��F����IU��!�jn�Uߦ�<n_���C�|-!���
�yit͠�iZ�s.��8�^ @�'b��j
��$hb�[s&��%l�*��[���l�w#��L#�7����>UmN�tp������H�������7ZtT�$�D��R���>����S�r����>A	�$�������ŏ˒
��1M1'|H�C��nð����+ �}9��t�^UI��#�I�>�����n�@,�cĒ�+��9:ܖ#���Sy2�f�����[�9�P��?0��*r�]�K���Ү?����--����CQ�[�R��ي3K�M}��趓=�Z�{ �Y�[��g�X��'�g]�ltK�y�]GR���[�	gea$��ʜ�;�/�;C�t��=�s@��KO"�����*|�]D7	C�PJ�����y)`z�^��G~��5�@�|-fś����cHXM���^�/j�lX%���I�/ЈK�R��	BC~*ߩʵhQɏe���=����0���!�<\�26��fS�u�� Q�1����[ޤ52�W�{�p�I��J#N�$�.7%���d��1(��z��9�V�|� ���.��E�$�{�H��AL���W,=���,�Fq���?�*�����4k�'��5���	0	�ǝmEL9j#�O�����i|��Њ����G�ҧ����߁�F���G_�(�0"�+��� h��ko�zv������,�ʻɽ]�� >*�7�{!��mLq�	�������-z�u���L79@�̼�'��8�9X哻�#���8N�@�j��Na
�/���*}����J�M��ʆ�܂ �}�֣��q�)Ҝ��3��dc.��(�-�7�����\��ą�Mu�䒥��XH�@l�]����E�z(��g`��Tu�)`������rx�n�ԝ���R-����6L�����`�Dܾ�0M�w�B�N�>E[���oΊ�T���DI��NO�|����>�D�����:P���82���`�}_Y'_[�R�����d\��D�XRzh˜W~?9����h7b�˪�T�:��|NO��r<�X�ʶ�3HD��|]�l�骼I��÷8�'I^�T�B���@�8�d+z/��x�Bi Sқ�Z�FL�@���<��������<��?z$D..{=���Y=��Y=�9N�~0��qkUg}h�M�:��mH�ć��ʊB�tn�ˤ�d�ks�s��J
?���W�$��u�U��:��kr5Y�ӥ)#���`|���('�:�h��������ke���W2�+P�r}I��3u|�du�]0q��n����U��J�C-_8rR��*�B{p#YzQ�(VV�1�7u������G}��mOF��C��%hh�!Ǔ��8�e�~��NMj�(cXF��B�(v쀒�N�a>\� *�뙛A3y�e lu�����9�4/�o���Sh�Y3�Xr�͠s�B�Er>m�j�s�4F=�O  ����j`6sc���P?�E�/�9�RҚX"P�9��c���(��I�����=�#�R�j���'0#���xQ�����Op����o��NAt�ڔ�2��n���5�&��9>Di�=*�۠HV~tz�V�`>�ؓh2u��8�	q�O�l}���Մ"�ʼ2�s�z�we��`��	���CP�GK��i��mPQ�tLt��@n���D/��w���Eig��[�L���o�X��*5��ݤ��� gW9yk��['-�mGV�����&��R�,�T���h�Sߊ��Gmc"���>�"�9m4�K�H01qO�Y�r}���\V	\�"���}�|z��VpD&������B
@�V�h�u�p��YUV��i�	c�� �ň�s����m3�V^���eؾ9:�\"
�'���t[�9B�ڑ���Ū|��3�չ)��O}F��p�/���h���8җ����1�
Ŕ@A�8���ūzZX�/bA�`g�	������*%��h=Ծ��cE��VQ��!~�g��Ȝ���D�/XpڸB��b���Nc�q¡��s�p�" X�����Cy��k�ʻՋ������#���7����[�k[�!�{Я��h� �V�^�;�����e�́��T}�xi����X�n����w:Cp��1ͫω�l�AFP���l�]{~�$�`�p�N�D�M����ҤV'.���!~-�ګ�@U%0�ղb�T��P�T����$ϒk��|	���Yw�����JS4��e�	�,Kq��áQV_��7���ݜ���L��8�#��TꌄL���NI3P��k�*)܍Z��^"���{�L���5�ʡz[�nK��Z��-?a�n}	>(lWj��E�U�.%�c�r�6Ǥ���ï�k�R�&�#X�b>��|���	w3F�;ᓿ�T�d�T����@������WC���7a��a��?�O��r�Q�ՓgU�ȍĖ�7�H;�X���&i	�yG�ҺPx��~�� �b՘dW��(�����h�w2��`�]s�͝��9P�ЪH�X9
�
�<���M��_.�����b㧓^KI���on�2�KrN�n�G�}���y���?(��'($;�c�9Z}H%l8ߕ�2'���j���]����d�w��v�v�#�z3��8���a1��k��l��$4%�������X�ѩl�J�%hWF&���똥��<� ,�P�d��U�[��_:n��r]7M)�r��c�y�2��q	�2�x�d/�纸�h "�R{��W@�nf6��+��8q"��;��V�(�1��,�`/o�7��	1��/I�(���#w�F^@�m28��q�!��\i�q����eN+��!G�{�]��N೟kr�G�,�cq��KFٶ�~�m��'�X!�P��J�cj���5N����$�>Πj�V����C"G +\���V�ܣ���.~�4�W[��qQ�|��&�UJ^+��b��?,ЇՔ���u�z.G݈���j�7�Y)����Ǉ�uyH�Z���/`�q�\x`����.�с���JJ��<�����ǑK�	���{������W35�e[���MZ�>�[�.q$�Ǧ�֙�.$ÄE�_��VUJa��X[+CO�V]?e4����� 40��)�"?����������Ʌ�f��T�� ��w[<E�C['s���dfUq�<£K,��۬.�,�<Y0s�su;�֓�+IZ�iHg�'K�%#jA��[����M�m�x���eM_\Q촴��E�Y �-J��bӇ7[ݜ�jr���'"�)W���u�u�w?ĝV]<��$D�����g�t�'~ż�g�/Q���N�u>�?�h�EK}��ŕ�m^�~/�Vf�XM�1�^��k�|"��'w0��9��!����~���5�n[�Ğ����d3_���:��=W�6��%$�q^���xd�s�� �na�nY#>�Mz6���O�ѿ�p�Jy���CW'�be�z����0����a�Z��O=c���H-�/��@��0����� ��5�����[���K�\���yr���k2���g ��o�KڪM<���N��q��w�x�-�k����1��J���@lg�֫ }�N:�Uԩ����;�}�P�
!BZ_�"��2�����G�Ck��@�{���L�övOG����s��t5�/��en���ɹ��h�<u��p�q��[���`�S��gm�0!�� \!���`��Е�U�l?o�y�ԅ�!������T�s}�@9
ǅ�P�l}���&�Y�#�X�q츬�}�"r���^7��P��������ؗ�D("�� ��>��G'�1pʒ�[�{�+Hj��=?�+�P�h�;f0$��2��	����dH�@|�B�w3����M���垎��k������{� )�=|���FUW��L�Wzt��6�Zg۵Ɉ���!j��������b�e��-��nMH��-������x���E���'���jύ�¸���EO\�=1��03�l}_�
[}x4��a	&l���h_����o	�79,5��痵���/��x�MU�N�%EȔy���	��p��)ilu�������O%v��k5gwj#�]4~��t�.X���-�yCZ�E'=u�=��P�DxVh?���U�z���^A ͍��X�~*�W,~�_Q��;Ə��N�qxK`,�s��Ѫ���'Q6���m��o� �W�CCۑ�����b�pW�AX���&Vո=��ڜa&_�c�pTI�[��E�TwAo	���&���wئ/4ϳi�"//��P+�2%C��W3<'1��%���I/��v鲪%&���z�y�<;ϻ�x��?�g�A>�@F�����h^"��,�r�c�ݸ�xA��!��t����j�89+밫����l�_�X$Y��"x�USC�aQ�}�����iL�Ar����kgX������F�Ql":3bL����x�oRs��=��bJwl�L��!OP��=h�/N��̈́�L�4��Ѫ��0����@�5��[8����"MJ��^��Pg�ʨ�z�ސ���Mg���9lG�Ez��(�ĵ(���ɮ{���C�SƓdP�M)���H^v��,��:q��r���O1�<pr�Y�K˚깼�33�"��x��V9A0��ŋ>��Ӭ7��胝X-��4=���]@��,~x�~y�!��掜�Sܘ2:�oy�ֳ�`o� 9�ҧ��y�K����p�N� H`�{��m��g����Td�G�=�F�Y��OF����m
��NL��6���F"���2 ��rK��?���z4o��Zzj����J�=��f�W0��~��9 G�7�M�c�R�0_�����,�vH�w�� \~�ʝP+	�����o֜wu��t����?˧,3�T���[�[V5����Z��۩{%�_�1��r���%�� d#���!���8#�@���g�!�D�:�܏j�%OZt�W�#�����ƅ�v�g�0���⫈xƫ�!�rG�V}߮�o��u$~q���±��B����h�uG�e�ЫQ9�`��Y<¡�K��4L��]^tP�����*
�}$�2	"e��ʉ}v݉���Q����z�V\�b�tvN�XVo  צp����8UQ&��`Ϧ���Zu���N�R�T�쌔d�Ia�:�'s���M��q�Qh�y^�0Z{�Yh�IΒ�����$nH����u��EG��ۆoZ��i&�D)Gm?Z��UT����M��@e�r�{��`�`���"	-,
��&�'^# iFh��;i�]O��B��Ѧ���3�{�৞o xOr�3P��Sŭ�f�H#:��d�j1!�9��8L����/�����R�c���s���+�}�b�������GV�ql�Yn�Iܩ�Zz�kg���/�Ͳj��/I��ǭ��xč��g1'okb����u{+?�c��>���P'���w�T�̶��-N��k����7��k±W!r�פ`Ca-�m�7�Z A@]a���"%	6p����$�BD����~J��Fg3������?�ϲl@[\��Dr������z��������k�jZG�>����m�������ɷO)�D<Q��_X��A���C%�["Ȱ��a�1�� ���1�0O�M�@�v�V�^�5��F:)3'���.��<YBB�kX�}�v���,�/�EwRic���l�쥋��iÑ��ĩWjl�S�Q��R�E^��y��{w�*S�iu&���g���~���Q�#�Qط����I���~�SUQq�gSa����a�ouh�qX���V��	�*��r
���X9o_=*�C�}��|�����o��X���Ol�� k3=�љ񒦚�G��X�]�[����Y�Z� �ڰ���v�D\.��5	G��fJ������c*�tTE�&<�d]p ��47��!t?�
?$1dj���H����FE?U3�ľ��A��xy���N�r��J֦�&(�}
t�#�,��N�Z��o�Eq��xMj���Ec d���/ʁ�f�nutE2Nb@a-5٧jmFR��z^+5��jw���.ë��;�m1Sp�[�m,��a�z"�W.o
*̿ �D�p�Τkh�z�'jPoxn���֜J�����3E2�R�Dkj�(-GO�ۣ��7P|9ۄhf��]lX��T�rJ�3���ͱ֢n�[8%ڬFj+�����'T��!YỦJC0�$��?ꁤwh|���HαɁ��������2xڭo�@K�U19h�����?�*A@��_���ry�*��y�����Cp���0�b��a{҄�`X�r��m	���>��_0
��<�Vt?3��4o)����dy"��Ʋz�5s#+�O�S�%M��7-��Ac a�b_��%�=�Y/l7f�,*�p�$�0�HV�
�(�8�yj���3��K)h>9�O�:diC�lK���L-�����81H,�����v;��3�_��~����h�C��G2�?���tk��#�n�&d�h=T���_��>4��v�lQ�1�u�ާe�!��aR.�d�4ั�-�BzM�h]��^�6_T��:標��#�[�l��L��	L7Q,�o����V�!������K����\t]"/p`�;c��j�+Z9#3�b��2��XO�������_�G��_KW�,d[΋�|��p���(�4��[��KK����4��&V�P��(�q��En���4������O�B8��V��YKP��܁�z;E����0�ߞx��+d�G�=�b�����U�
�,�6�K7nv���t�0�7#����4`��q�:=���gzW��MX��s�k�f�D��z�����w���~�g����6n�0��N2O�h0��bvVX��A��I�Z_^U��i�����@7�5��j�%\n���[~	� ݈�w���^T�]�%`�ڡw;�l25�O�̗������C�	�����+ h`������GV�q%������d���|Tt�M7ӡ� �G�ڕrr̈?�\�b�`�W^`�#��OH��Z��.V���5�Z�Y���*[�i�v��S�����Fo�F���:H<�����^L���zM>ط�d�4~ >�Z��r5\��'���~��I[�d��Ru���=Dޤ6�������i�]3�]��~�b$�P��h�-���	č�+NU��«�e�ܚql1�t4�3��W\���rS�	�R����1�R�r�����x}:`�[���c�.Z������݀'�1��p�U�^�<zLT.�B��F<���6��j����WS;�$x߀V����g�9!���%�G�%��?�s�W�8��w�W	�d��Μr�+I�)�qh�S�Օ7zzZO���wZ�7k����p�D�$ő��ˤ���)"gf�SR�x��C�}iއ��H>JwT��_���V����:�l�"��N�>��4Aӄn_Z�ˇ�Vb)�w
'�F�/�"����)�"z�
�Z�T�B
@M���5'Ӌ�M�نɏ�)ʀ�-Rf�S�֢(ҳC��;P��Ǜ��pR4�rl�-5�\! ��n�X 0����7�RV'�h�+��0� 3f)�1ym�Jj4`���+��:��_K��4-�ے�#��B0T��[2k#�Q�����"�g-�gI��ɝQ���Uv��qx�E1h��i�b��CPO�	����v^�&�,��xܗn��T{��}����2�S#��1p����!n+�`@����]�R'M���|�ɲ��7��g:���p0I98.b��M�7�X��\��0!1����Wm����f��쫆���
�(�Ʈ0�w/Fv�^mLͻY���_ç[6�4�@��I��b��ǡ�L����^G���_�3i֠�8ݱ]� ����Y&�o('�����<�6ó��q�v�N��CFag�F���ǫ"\�sL4�~������ڔ���R�niED����C�?$��$�q[hR��:�}�U/c��t/�
�%s�k��e�V8y �3M�&���V;(V�@[nD�}��ދ��N?��C�۟�;9r!#,�qW����E�.���5���N���e�4�����ar�cp+#ϐW���{���g�%h~�Y�8�����}���uD���<V� ���w;L��jf��v*Rɉ�^R��I�d�����|�a�]�ņP��������j�|��@|A�j��-���kj{;�C�b�2x
]��`G5���)t%C+fc�]��P�.��ס@}� �%=ڹ�Un�����/G]tM%���~�����0H����rz��Ԡ�@ݪ�A�Ҷa�3$qܖ�A��,hI}�u�'U��.ZJ�2�:�H�g�6gY�M�7�#�G��w�&4��p��L��z}�i�\
�߲�m��f���(q�q&|6�E��u�uo�(
���pyU r
�_:*�(�P���\��'�?[�u�P7�5���e�I�Cb<n6ȤRr�` �az�l��L�r��m�����>� �	��Y����`�?����
�b�>���'��M�_]�a�f,�DuE�eu2��`��V�M7�6~Z=<�9�|i�Π{��Цr<ai�-����_9��T�5�`���u��e![1 ��YS�zR�&�����&�O覮9�����+ �8����,��l*Oɭ�<4�A��t������*�Ï!�"��8��P��g����4�9��d��#,��+���gs��5)].�5�D(g��|�e�氶(��������R�@2�4X+jֵ�xb�d��� w�'p�ڀ�h�l'�,����Q���=����]g��&������z��d���啂AM��p�R´���w� ��/K����,:ֻB�`���SkJ��-���,I�O��s��OK��%��#gT yǳ���Σ:��1}�%�Q8,��E��H���t]5;og$U܉"dP�K>d��(�^�;���ƿ�	!P3,(�K�_�T=W�2�0�����*�1'LΫ�a8 ���SJ0��R���8�s΃T Zv��T�yL�R筄hBa���W����Fʓ�i�ŤQp�˦�Y�R�ϡ{\�jOPK��Dg���q���$����BNѥT�����A!E+5G������+�]��u���>tu�x����G�v���+�r�9Q���i�;�T�~�.ɻ�R�� +^�h�TT�L躱�[����?z�"�&{��+uwi�^a�|�;�,i��aX���n��@_��b�)V�ʵ��r�͋!Rr�p.,���xX\����Vx�$0Ң���w(�V��pǙ� (Q��b.֬S��09�Q�� &cK�����g.
P8�2md���#��G�����)U�L������O5o
�����Z�Sj�W���b�I�i"h��-\̬m�u���)���N`bgmH�w��Y(>�|{=H?A��:U2b�³�W�b"V����ޤf_ԥ+��P ��w��!�c�6��Ylw�λ�W��Z�����u����ߖ#��K�j�kbJ��}�c�7��|l���	��'�
�kcgAzV�THm7^��	�ѸWӹ~�� O.���~(��!Eȴ��JR��ָщc�L���,.D�eu��GS�j04V�(\��O�RRif�kĔ�(�;R�ǡg�S$�� ����Q��uH�Q́[��ݸL����㗻FM=��-�eMVI���nO��,� ���׺"�N;�)��;���{�V�rF�K�.P����V�wq�zt�6���2�������n���[��#?��1tI6漀o�v=�dA��RF3��؛Ŵ"�A=��@�Й�Mט���:��{�9k����	W4�ͦ�f���/RU5xm~eZmȳ��h��ġ�#�qA���6l��BU�^��� O���5��ͻ-��&��{:�hx7jݬ�YU�M�>�$�1j�K���g�Ԟ��v��N1��:j�w@�M r7Z6]p(HC���R�җT�@�BF����K�ŕ�_�Zb�)Ǐ��Fr�#�}�[�w,ĩ�#�feŋL\�8��w�v�a�I�U�}M��P>+��=Gj4�IU��'��g���z�V�Ř�(�c,��@p�����D^�~�}%\'#�Bt\����}j���[��t�6E�j<��e���?�� s�*l-<x��8S���ʌ'����ױ��g�9�{�����AizT��k����"$�I9ϼ~hR��H*F��P/���_�&Sj�FW�5Ò�%���8���s�˯�z�(�g_x�|�*�J�`ʡ��b¶����7F<E��h�"-�K�*����hL@.��������4*Q��s���	�pY�|�L������c��0� B���񸣸��ĊF.�<v�_�_����>��H#Ѽ�kgs��8yY����gr4g���sO����]�d0{CV���m����a�3P�&҉�����K*{+����)���`�T���E�ti�m�\���)��x{z�7Y=��pz����[�+'U4��.�'��,X�B���$��x����.��7"�1�6�Et��wX(<v�Y�E�=�h[��Jv�w�|��4��#�̋�`"�\��sѾ('��HJ��ri���!|l�
e���_}�.\��4$�)8�;[Nf넒1���"�w?ۓ�h\��4D��ݢ��:^�,�u}_�3�B�� '�V�en�yu�5�픾ُ�t��s�4�,@��Hi(���:��P|�G�洝����I�ط�������~]n��<:���bx�����^G�G5/���|F���Q�g������]r"��U�;�� m�$Ax�~�o�|�`=ŝ���mY�G���$ȸ�L��mA�p���9�_g�p����=Ig`O�pu�.<�����:��S>���	��9闦�f�/��>N�k��_轞��������=��oK΄���b�,,lX*����Z+19A����=���˾�K��$�"AE�]��Jl�A!�4hP����>�
�S~1r��o (F���Y�"��O�-~�A '\�j���|��a�C? ���%�o����:���,Aw��J�îR�=�\rjc��w�{�"��A�\���"�Wu�ucm���6�d٢���*s��h���n�.�5��-��;O�A<�����R)~u$Z�:��9���h��z��6A��F�P�Ne���A���vHF�.�� n�2��2�p���.ܴ������H�p%�v䂝Γ���;���n�� � �_ցx3h�Tyz�0O���v��/)z�I���QeLdj?���{:���2���\�}an���LV��WV�tq������������ӆ���Gsx�.����( ��ǻ�tŹ��8acd�@n:c!����?���V�<ħ���k�ZQ��O���d�D��Qk\ �@�S�9�+jsd?�n��vu����bV�l� }X��0��hi��Z�NMsICb��`��b�G�G�=�x�b�"s�lϡ�eq#"���K,�2Y�f^�P+k��` ���3��nv��l4(�%%�Q����N�)�	[��G�h�<4޺pU�-�AAu!�����c"��U*?��E���J専Is5)��YH�4 �h���*}Ы��ې_�Ҍ3X�в&pD��k������S^&g��+�+�}ںƌ�������d��3.8N	��%G�/��Q��5�8Ǔ_�Y���q`g��m#��*�\i��4f ��������� P�"�)�#���N�|��d(0�;"ޝg��y������fȒ|@���	0@#w$K'�F�%׋�+O���R����k�gS5| l<\<�HU����	Y*��1}KO���xO6v[�����l�pR� ���j�HL��1�����b/xeW�X�7�Ȯ�'��
�𔠄Le���+�º����W~{-��|�G�_})D:��~f�F�X�����?ϻ���)�s������z�h�oj6L]A��w��n	���ss��h��&(�a���vQ�;Cy7�^3����*\��F�6ĺ�d&� ��������\ݙ0�1b\����J!o�w�(���Fhr��@����P�$�?x���op�Z��a(8����}�E��z!�q�@ _Y�tn�w�ʢ�ݒEC�TG�;
و�&�t�?x_�i�˲x��_N�N����~">̽�S�)AQ�=PN}2b���i������v��14���	��Q4�A����	x�x2ld� �{�`��?����;���f/X6Nv7`���.���aj&C�1%6o�V|*Z�k�.�K:(j�	���zB�]��&6/KB@T�U�\VB�Q���w�M�!E���L��#i��~���^s!��k���@Z�
�Z���F!���Y�D��ɛ�q�
�Іy�H)1-i�:��Z��c����U�����76�t�U�5�.�#q��:�,"��V����Ѐ�}�������t���M;���EYI���.q�r����ko|W��9^��"�J��[*���DqmV���I}��0k���(,�=�؆P��f�N������˱���)��l�D���7� �t��k�p���e闔�r9��2�a(V7<�)`S����>��9�*uqVAS��חdXu rG��y���za�������j��mxTw���/��us9�Y����ySե��� Z������-��'�FwE������n�&<! nOWj+����&~0��"W-�6�4��O��&X�ȏ��UD�f2]ω����A<���u.a ���-Y	��g~�H;�k�6���(4�8��8iq_�S���=���ؖ�PF��1�	*�j������R]�;�'���3S���	��6D7�Hd�2��NyroG("t��|lsIOzA����MDb�lޥݲ0�5���3۶B�j���ZK���f��߷b֑��S���)Y�2���w�U�Si������Ed���ܮ�Y�-(���`ɻ_i<���Y��6V���=�8��@l��b�M$�'Io�ly7<N��[�F��(緪�I���eٳ�#��37>�m^��ڧb|�`Q��;�#H�;�S�J<?d���B�C�2T�G8���U(c@2�ͮ����TU�� ,U�wgxA�bӯ}�ϊ�����O�4�A�
#B腟`�i�q�����W��]�A��9�w/)�؞��V��K�!z�)��ݏ���(�x OOaf��A�5_�?��rE�e�yu�NX@���]���w,�\!��m�|��+�|�VTRFҐ̫��7�u1��su�hUp�2�F��^_2��J�p�~�.��5��L0�}kR�'[u,G�3��ߏ�a�sRN�����?�zm����rw,�r��fQ�OM�o&��q��U%dV��q�C�7��c_�t`[ٛ���ä��Y�'t'�u�)��0y��Y�����m������ͧ������.���sStPg��Yj1�v}j�KL�X�^q{5��4_�[�n7��h�(�2P	¸���E������W2H���e�
����>�7�l��&#r���cC��~$�R��]C�R[��8���i+�����&,�?+Fy_�"s�9��c�;g�)S�6[�;Y�&i����vh�ˡ�-X!�;����,�
,!�"�	�FpJ�Mz��_�J�G4���s�ߐ���5�&�DjQѾӱ��}�%	��p�g�ѩ-���q\N�C����+3�Ea�rp!\����Z���þ�����5�)و���rH2N���q���1��[bH��R���r����������HW#������O<�O�"�}�\V2(�IrA(�	�O���uk��,Q�R[������(l���{����Qۋ�v��ź�,�~��7�I�+_X�]���� ��+��y�/B��r0�C��?L\�W��3�Cq��?���8��9�s��Z�GW���W���_ԗ�XIX��d����X��2H��{��&��b�[Ыk=�ʀ��؉|�X��n��K���+b��Nn�����YFv�ܴdRrɱ�+����f�=����F���Q�oR��{t0�h��D3��ďSև��%�m'��e���n=J�OH?��e��͡�R����^r!�kG�j� ZT�ގ�]R�R�h1����^��/6f4�Jԋ}H_�
ƶ85�uS�D��h�K�g�ʍm ��u�W��eU��^���f�^a����V�K�lP���Ҳ��<�t�Q9�P\W8f�<�y5V�cI;�;�ӠO��k.���%bp�	�ؙB��Z�|��c�U��@����'�wQI�S蛗�̏�f��g�
�����j������k�\-�7�q�ؚ��0�4���@�E<�_Ptcg)�r�o�k�Xg�~���-��d_kVw�Lj#;f/�.��g����Y�X��S�n�x��$zM&�D�K`ȧ�D�$Uj"בa��!��~��cH,�mU���&L��p � R�9G�J�G�!4��m��v~�����]n��9x3NÆW����*Nº'=v< �~1��&�����9��Qw3�X %����\���\�vb�U2A�x�u��7!��U_R;v'��<䊑d���{��Ϫ�[]A]�Fl��v	� +�Q�����p�-Fd��RtC��&64����P�a=��Q���$z����[�+3�$�e�4(,cf^y&�NSZd���h������Y��kv��_�~����>F��>����̷�LE��-uM�
hR�a8c��/��Ĺ�p��/h�b~,7ǩ��Ya�����Y�n��	�;;�TR$�t�K��
c�L�8��o���Go�TF�NuB��"��jv
 1�,��#�]1�;���N�dz�aZe�N%";X!���ⓞg�j�<�r��7 !F����\�F�9���?by�ᜧ;9,F��ۗ�`(�������H�ׁ�b~��o2W�o�����}
��~���%�P��Ԧ���r
���"��i�8E/�Q:��.��J�D&5���a��Sp8�`qlX��gi����{���>��
R��|��a@���
�V\��R��g�u�~�se٩w`��ޮ�7� C��`�8e5���0�%���QD����KOd�p�GG����-�%��r�{�u�(�
?�3hd=�?�K���|yTE�=�㫇��?%�L/ŀB��9�G	�FbެL�6�h+�,4X�!1!�ԙ4������*��XÙ��0����-^a�3+N���+1w�|A-FE��I�Of���P,���#a�%�Lݰ�w�Y@�~�SK�B�L�����Cʕ.kv6�Of5����qLH3��5����=�f�fu\���8B$�� YT0s�-����u���8����ϕ���
!��.`^�TR�+tL\�<���K�������Q���,�$�ƻ�λ�ʒ�^~�ݣ��JS���!�Yi�B��|W�|�){�+��a��w�:�pݳy�L����*�$�zٗO/M�ʤ#�-��Vɪ<u���$���r#�o�TKG�WU9�,����qc"�o'/��:�/��x���/��X�a���Scl�OՏ@�l����[Q�눧^*���"8�:��GR���H�=��Iҡ|����H����^G�aZ/�[p�Ʀ��b�K��.��Z=b���	�m��+O�=0:%��Ѡ4��@�	�[V�OW~��!���a���`�?�͎ҿ�"���?�� ^l���_�o����f��Cn��`fw�&�y��G��3nҪ�۾��"��	�p�;YP��;1K7�Z�6PUh9�����Y?;��F=PH�[�]Qp��b�m����B�i���)�د���읙OҚ 8�d8Pr7h�Ǒ�?�g;	�)&^k(z�u!�O~�Xu�[�7D]_�`&/dvU����n�0���ҝ�>�]~Z�C�[���A�{�	�D�f��X����e@�$�ģs�!Eܫ������:�pw|��p�1����CUn�>;F�<�a�(p��\�&ՠB��Ra�D��#�qOv��0�%��k<����}�Z����Z��羽���X�5F%�5�	�.oA��2��zfr�cl?��9�\�\�c{H�e]qA|=7�y��� �?�3�'j9�S[M}��YD�D2k�?�s�j�nj/r#>[�OA���3���,��m��O@�av�h>X`<��ܿg�u���ZyK��1���3�a/��]���A{�Y7��{��{��V���X�����{���R�4�e��а�z���6a@)t�Zb��-J�3���O��A�̩{{Xv�q�9Tl��ξ�����M�\P~��m�8��d���F{J��
rr#)>	��|!�B��Twۯ-"M���C(ۀHZ2�^��a�h6g,�����i}��M{?�ج�5���͵�����
���o����al_�K�� x/[g\�Y���(����St��_������<T�����͚؁~--����ϔ?�$M4C��|jȺ4.�uT�m{{��XX����@�T�$M]�g	�����L|���z���R%ٕg��U��\��}M��O��l�N�Yi�������=B��":q��h_p�"���㕸D5=?f���3���uD�����Yk������b�b4��vbsZ�����k����!�fç�qM�ښ34�!�U*[�W��^�s[|�p���J����ퟅ�O�V�_��0u
��~%���虝�"�s���~S�(Dq�&���,x��S���������]LWT��kcY(��2��n3w�#��i��l8{ݥfK�P@,~��lՂ�C#*�P��:	.sfG�%����|�"X�[����nP�b��o�,X���-��L��*�X(?o�T����s�׭+͇J�^��zV�=��~G�-��C�qGL3+��oJ�d:���0a���t�wu�-:N�I!H�O4���%X�O�L���i���2��w̱�H�-'��ox>��R�뛩�y�lv��&et��x+^~ٓ�M�щvK,<�l: 1���B
)��	����П/t��¿��^<���fƳ8Y�[�JK�Lc.��:b�P����;�@��9[dL�N���O�4�Ԕ2HB���y%���n��φ��
jS�p��)�Ơ�w{�c�'9��1��V�tY��l<&�p����c�|=��}��5����*sgpty~L��y���듒���d5��^p u��l�f�Q� �W�a�F���0�b�ĸ�gN��
�����i�42���a�H����'jO�h� Cژ�DޠG��?�V. �­X��nG�N���wY�:�p"y�(�r��~W��ۏ�ZDeY�Î�r�8�}��U(��an�Z��{כbi�w_�Ti�F_�12<���(���W����gY��/a���b��zM�(j�:����7����E#E�:q�#�n��ʎb�M�P����?����H�6�.0�&��Ԕ�+E�3O��})=��u%ɫ����6��Ҟ�f�Il��G���GU
k���"�hr����2�F:nB(5ߴ) մM�A<�UFys�v'���{����- ,���ƼykU�~V�j@�11Sw�|ʗ�x���u��8�6�8~�~M��[K��?���}��R��[̜�ƕ�j'��Ϋ/�yn�|L�@ݱ����I���5�X����풿�,#��q����F��%j���l 8�(�-E�5�C��YTMc���o�wan�k�l���P�f�,���)wW�1J��|U�'�����Z
��h �OtT؝�u��3� ��D�?5���������}A�ET�]�<��L�:]��I@�U�ڕ
{�u$I[�	�M���?��ms/�6�i���J6{�dg5,~d>��s�Dϕ伞���j�ƶ���g�^���c3�s���$��pvM��fQ����Zs��I�����L��~�&ɾ����Q�6��yՠ��p!2Q�MƦ7��j���M�� 9��e�j�Y+w^.�����y�H/�G�9W�$w�c���F�j�j7C���>4�.����1�"2 �)�OXΣ'��1��pگ�/�CQc�J�m�4��l1Yy�_m~�G�a6��g�
-�`�򈺖~��h>V��h����/��2al�_B����}Q�ft:T+tC�\��4�ƃ��L�@���*x���� -�2���=C�έc�+��ߐ�$��'�%��\�>��M1|ϴ�m��Ԓ�[L/،ds:�Ú�,���V@�w����}-hp��tZ�|�b��-_�!K&�A�>��y�[����N���%�"�;�N����B���P����Eq��d+}�O���T �v�:�O��+�'�$���� (������2�~�[�����B��
Dd����?�hZ��]��FV�Gu[<�l
�A�>��aX�<��tQ�+j��� ~알�2 %
y� X4L����������y x��VT��o��K;��	M�^5��^%�^��oM�m��y�xu-�B� *������-�����<�y�&.@.��w��f.�Z��	����H?B?��B\�#�Z}�FR!�w��S��*���j{>��
�A�һ��l>h���L^��V�_�����ep����R�C�.Xo1~���j�p���E���	��7��>&�h�gi^�WG��6������/j(y���~/W�N���	�W�h��7e�u����+T�vކ~����wBF�0cm�|�!PH7%�%�p�qpg�}�\pؒu��%��i��i����P�?QH� DD��J�$a5� �jZ��vy�9Vh�Rܝ������E���n�0��_���F�μ�v�~Um������4�e0�\b^2ڀ"٭�Z�M� @vW%��Yi�]���m�(�k
L�ɲ"�Ԙ�O�'��ᓄ (;Z>:�S$P�5���j9�-9��Xt�mt�MJ�|�j�8�=��z=����ݻ�A���ۃp��?�uv�g��@�X9�$�j�U0��� [�Pi�~b��z�._�#܍{*��R����'z�;�Ԉ�/&�k�q��[a�kClY��,(97gedɓW'⽒�.Ը9Hu!q ��jQ��e$��C� Lb*�Ŋ��ex��u��DB>R+پ�_��D ʃ�*�ܑC�/s��/kk����[�M�w:��5k��u�ɍ�.�p*s@[`~��_�e��T��Ɣ�j���g�ԩ������C��/ޢ3F��Jƍ�e��? 6�^F7����m_�Q���U��njU�z�dЕ7�O�#�ӥ��G�b��%+�Z�k�1���&�� ���V�]L�~}�p�B��KsF6�+��4_ʃ�2�{O��x�D	-����=p�x6�F���E��Z*E89%�s���C��(	߭��'ȳ7vY'�(+��e��7�5���D͸VyE�$�3�3�y�a�󘼍�K��L/�����/*y>v��P���:V���FB�E�g��c?5��ez�ig��+v�����jT�t�A�n�赧YDĩ1B=�ӣG'F	�D�.d�b�$�/ <��1��&;�rB��<S/�[[3�[��[���6R��y��}�t�6|��B����˟D;�o�7��c��\�>�֠P�E���T@ܣ�I?:\����RWSvN���ՠj���)�#/�!? Ƀ���]��fա��������#���丶#�����a?�����iK1H�#F�&ԧ_�% ;{2�T=�>�V����Y4Ne����+$�z���:�m���/1�"#0��m���?0v�h��Y�e��2S��f�<�Y��T��F�L�G.�I%:IV?�%?̏��z�/ܥl�l��h�^���v_��7�b�Bd��/�NM�J�x�R�a�,cֆ����G����𨝷#��ĎD��9-�Os?)$Th��QZ�99>\�Wy�:��j�Ǉ��>,����Gld��[Tƈ��S�a��,�K~;�>��ǌ�?��Ɋ+Ϡ�8�(^n�pZIe[ ��Ғw�3Vk����^ֺ��
���[�B�V���}�ۘ7.��8��[]���kZ\h7��iOڜ�i}���-S@��3*�i�"j��Ch܄��b���M�$$���}8������?_1ʜ�e2I/U��@z����&�D"�eF(��3�ނ�N�q����ϫr5��S��9e�I�CjA^�RW�.�f�p��/�7(��aQ�ۘ�1�$Q�͟�����^��{� �
��
�	��1��u��h������𙛞�5����o"	8 ���pb����t*���:��-\?�HEV���d�@�g���lܗ;�{��H�����M��%v.i���@yp�o�H���͒�<��E��B& ���sj�sF���S��?�+pUs�c׎l�*��Ҫ!�d�Z��A��a 6.����j.�=���!n�˷%�G���$� �V��2�/M�
��|�
�H}�%����r15�*������ﷶ�}����:�2�(��h�1p�e�Z��&عOr��3�w���Ջ���Y=?��'m*K�,5�L�g�$��,�a$�pM�v��/�U�ze��g�����ɨQ�=�H���'R52�Gi|�O��:��X?\�G�_\�}�
Z�f0��`����Y��3J�,Д��<���u�o���;���������Ĕ�u_�a�]y�������|����jVT���Xx�����rZ�T2L=��Է����ƭ�Vfn�;�*�8J��b�KU����қ��ӑj�0i+�mЏ��ט.Ԧ��Lx���El���h˯�����^���M?}���|������k0/�O,),=!�7�OE�Om+ڔ����Q���(�W��&g;g��&�6�4��U(�u��bZ�J^���b��)�~dy�ʔ��j���E�p��~�χ���\)ϱ��(K|����5i��+�8���_Sպ@��P��m��$яǶL1#2�8�����y.���w-�r;�*OZZ�$�}���-���ɝ%L#y(���&�N�����$���{�|�!��KRܗQ���'�$LW�����#�bC$&,fu]��,i�ۨ�.w���_��1�<痶��q-�m�@����g��z�<01��g\,��_}�a�+m)l/՟E/2̬8�\��Ҳ�����JB��q�K@G�A�C���9�)���9��+�O�Z�n3x�s1�ouy�5���n�b	jV�':�1���"˶�3*/Lw��O��%�Z9�c=��K��2�:��HAH�?�k�����Qh倄�{'��xs�3@ �eƣ,3����I���Q�U^xw.?��8�dcI:䭗nt �{Z�p�7�M��'�Q�L ��b��Q�Y�\�q9����>&� �|��#�@U��r��T1FT�(��k�d��D�Q.���n+_䉡�����KL��O�D�w�!�l���i#�v�X�ޯs���D�p����R���l�����Ѱ#C�}�D.J��ӔoA�:U�b�r�M+5��9��'2O[�`�#�L��sA3E����3{:����[�i�4��}��<�/#X.L���8۔��EAs.d��;\�T(�� NP,�3���JR�X��rTY�z���|/�kr(����XA���k�c�Ok��G�����lŋ$�,��a&$��@�8�;��;p�-�]V��X9��G�!%M��=z"� �,�i82fL���[.M�T��������4Un��ewyu�B]��\�AƂ	�[���a֚�4_L�3��sX����Q�Φz�]�����a�j�_�1�Qw$y@T ��P���hi�ܪ���Q�XB$���|$~Trf-h��}���ǌ�w�i�|�I����R=Aa�s&���P���U��v�+VX�[d������X��P*��[
��F�j�R�1c�k��$VN�O��~�T4�����-Z./�"�6�.f�l��AR�[�>��Z��'=*�S��@�U-���r"���9��<��ZX�x��=^���{������p�?@=��BvԽ��c���	� XJk����t2�Ж���P`e
�b�OB���^��?%F�������`�L�^l�I�|�a.�kvϙl覇�zr�~�Ha�Y�l|5��A3q���9I`4g/���;0-IbztNk�Ae�v��^x�N���E�,5kR�EI �$Sr�!���;���l�G@��|�e�[��č�����ҡ�C�ͭ�|7�z�Y�X�(��,��.k�eܳXH�\똟5�V~г����iM�eM�,���ⷾPW���#ݪŵaX��M
��0�{i��iB�rN^n�m|��~K?Egh
]�8��8/*IPƍy=�[����G�m�,A��uDf΅u�u�&�H�<gY��P�*�\+h�;M�aHp��'Ŷ��K�S8�|
[��HqS��S9B.dY�C3����>?�'��(u��G@%���.9��&���^)2�_&©�[��*U�ܗ�:V2-;�;��FZ��������*�xФJf:g���mr���! ����\��"���T�b5�L���^r�ծc���b��QG�S:���f��6; |�$_�6\~ef<~OP���5c򩚈�F�d�Ib�2�Z�̭����*{o��n+�,���{]��C�9��P�O�ȕr�����FA�T���\���6LLM	_�7�W��7蚷�⌌c	���Dg�,a�ǉ���I�XyUX?������Ǹ��UOj�4��t���SN��,��H��z����[�~P9�ل8���1���ȝ�nJ�s~��];,�֥��/�Wn��*���5\�@��S0|H0�K�*�t��J�2^(vY���y.SW�RAӐ*Qk���`�r�٭mF<]���1�S���u�"N�����X�mA,�RO��<$#��N�Z���im��^2�cc9�
%�L������.t|�s:�u�M�-�9@��scq��1��M��A�Ϸ��p��P���Ɋ�S�'���Qmu����7�K�5�Z��
�dA����f�'R6�5k�$~����|����Ćb$Ǌ�I�m&bPOm6�U��gDƷ	,0�	�&��4���`�b���-p֖hN� [����:��z+�\v8
���xl������0F��ϵOX�(Z��Ew[��K#g�����3�����ikP�.���lw\D�!��͒=�2Ke���� B/�7ۥI
����V���s���ٵ&}�D��"Ǿ��}o�U!�[nB	��VѬx���R��t�%����d�2U�F�R�H��}���PS�XE�x�"�_�N��Te��M���;�K~���!q��.�^�Ü7���Z}W(�z���^ !د���~�f2�&C}��`E��w/(%�8f�����a=$m�]�H`�ٚ���F{2u��G������b�����H��T��nZ��}[�'t|�>�&��d���f⋊�%�oN�",�,w�oQ�,�"a]�,4^�*G2������ϣ&
ñ����d�ֳ�x�J�V���P]Zmeڿmz8�y:`���(^b��I��&K*��sl��4;@�N&�G���8*ݧ`:׳l�Z�-�b�c���R����e�c)�m�ҝ^ ��A-?�Jd���>E�̽KK�9|o����Q�n��T��	�ן�`FE��<�7���i��zʄ��(H8]��Ib�Lv���_H��0��
��rz�ޭUP��4D��	vy"(�����d���� ;�i����4Eֲ9{D/��}O���0N����D�;f�ǵӺL|�~�Y&�?����T`x���R��x�����?1���������R�����D�3^�;:�F+��J�����
ט��,dj̎�KH�EANWZ'�Yá�%��P�cz���u�tS	��n>~��T�i4����.��'���%i�1�<��M��(���^����#V!�e{��*DwDJ��h9S#Ѐoܗ\�A���6�~�Sk|	O��^�#�P�)#0�]hg9G�׃��sg?�~3��k\�s�r�v����#ثV�h�ڇ��5���[�I�A�8�A4��^��hȧx!�s��
i;�z�k}������o]��L��_ �~Ư7����)�>�����XT��q:���bm�0��F�L^��x!�5��B��@�NmԺ�g��̜����d?'��h� �9qo)����Vc��S�$�/��|�h����js����BoB�%;����i){�W��w[�80a����i�����\C)�?F�|�h$����}i��n�թ����7@�o���] �
kF�����r�3��H��w�p�1~��iժV�Ì*iSw*����Ʉ��<�H@�81c�_�ȴ/��G��vT�u�n��AW[�7�W�JK��������o �Y%c���l�#Kˈ�'�먠)��Vm��}4�Z51⍶=ֹ,������	�j=A�g���o��U[S���Kms'_g��cF�BCzfJ�Ɔ��-&��O�a�yVŨӓ��H�
	H�/)R&B����ig�(3��֒�gm���x� �t�b�i[J䕳z�ҿ/�DL
�ݝ��TP[���5��\_R��N��Y�?��g��EN�ďWM���F��B;Z١�.Е�>7�	�`�$c)�+3�tY����]7��(s�6MH2n�|��W��Ы��H�M��5VS��6}����dE@~A"�"B]�(cw(F��غ�/ͤaǁ�Gg	Jw��gY*P"}H��s�*�x\;�X��Z���_ܚem�疵Vɤ��ؑE�Ʊ���2�$Ƣ�c�{�j�G�?��-��մ�`�V�0�+Up֊cl�\Q(a�i&�4��R�掁�d�;,7kqi�Ū&M(8(�����@��饠B�����X��*J����-��F�����z��@Gi���gEG*��Z�v/���Nu@��j&]�(�=\�Ƌu�C�x��`��LBi��Q}޺;��a5��%��E}�%"3����N�4C���.��K"�D'��Ą�8L�;[踕7�ڥV�?��C]�� =�1<x�[a��v��䵭 ���S���q�ʡ��˙:w=����Z1��u��[�pVJ8��N�r�L7�����U�Fvk"$��_�~�4���5�!�i���&cʉ�Q�����*B@�%H�r~M���Hz,���X�
�ӦYH���@�x.p�S0�+�����B��	Ȟ�r���Vc�eԍ���!ī�U��~i�L� ��2FB&E�y�S�yk\z�(n��{���\��|��&�+y�N������x��G?�~�	4ܘ�47d������Z�tL���[�d*ƾ��
F,C�	��nK��ޓߒX�F�Ց���䏤��t�XJeg`�rgd�"0߼)(u���@��7�*��C�D�y����յ�<X�DVb�0{4����L�&~���g�k\#v�ZN�#�=�t&&'Vr�!��{Ը�̉,(�@��R��.q�I�O��o��4y��#w�{e=z�f@��Fܰ�e'wGW�f@b�?����()�r�����9ߕ�
�̝ܱ���dX�pE�F�u�i�̇/�����*W���2=DY1�:�8�,s��)�.������O͈���:� ����B�%��ʹ$]_��}Cn���$�߮X������b���
/�L�4�G}KM������G����i:�v́!�S��ph�R���1.�A}��`o� :��U��iok7z�*f��Rr/'u� 'hӹ�+�m���Ʒ�x��cj0إ�L�H���ƒ���1���}Q��"{
G��(%#�f���(gw��#=ÎRB�˯]x��8n���r
�����"H���A�>h��)���?j��؆b:z�Z��iݠh��o�Ϸ�2�8{�����ўc$y��|<;R��o7�_��m�� \rC�u�Xaw��'F����_�����������˫CCЄ�ly����-թ����W����`���=f��/̚�Nī�W��MW���	���2�e�!F�k30!�J��v�U��+�Z��I�Q	p�K;�h$��%;�֠U!$��u�$�2�-v�,(�����Ѕ
?)�VvO��y?,��g��`ۉ�Q�Vw��~\L�YvA؁����ju�ˈF�~���Ɲp�f�I{����J��J�m�
:��{yJzT�5%Q���3c!P/���H��DT�]Is����>�c;{��</H���^�[������+`��F�F�6O�ۑ6m���𣈅�����\nzY�\H�0�2EP�:�5�5��Grߺ@,eL#�E.�"DN���L��rL�f�H�����0��yNv+�
���f�^X�Bq��:���?�)�%�K	�Rmg
�V+;r�e�:w�qc���10	ظ�;cI�ό�:���{r���akˈ�{�6뗸���RƤ���47�A*��(p���8�$�>v2[�/�Y�`��qb�d��n��4�C7Z��M3�<�:¯�&avέV�01�e�К��q�Z��^/�A�����P�]�����2y��j�4#)�X���Q����y�wҌ��C���
$��1Ԏ�qt��K�	 l�m�5Ec��T��	_ͼ�P'���\�=j���~AB�d+-�K98L�1�y�J`�`�J���O��o,���1�qv� ����R �b��M3�ǄO����ߚ]�/�E�sI�~��ǐ
,A���_<m����ը�}��j��Q�p�����U�s��~��UR-+'V�R�"��/hr.����1�'�����d��Ŗ���&|BY�W-�������mNs�fө�^,T[qh�pr�l���ZF\�.��R�F��`3`>52�\�f�f(���'R�ҷ� ȍ1�I7�鞩�r���f�%�2fXz��%g�u%�����Bm]��A���Nҁ�%���责�G=�(p��'��$C��d	�~��[X�=Gы��a��}e"�.�у�	Q�����?��Š��!7n&�J�� �c�Z�Mt,'_0�h��DyEccj���B����T�	xWPڵ"J��N	�e�zY���ƌ��"^����M��6O��~X���Hl
$γ`[��z�7��8�4��Xi��=d�SY�eW�>���Fj��u^�i	ĳ"�VHm� ��C�5�A�I�1iE��?�����1Ix����LaE����o!��/�pk��3���{�����7��xY{��W7�]��T���?6�ޘ�r��d��4���Qڃ�a�+�9Dq�(�Z�#�#��~@wK�Gg��I5r�	\���w��Ք<Bx'���˃<�a���J4��MÃ����%�1�9�gj��O�����U=�fBO�>w����J��`��ӂ�K1x0�[�"avh��g�0�ԭLT��]�	Zž5�a��Ӫ�M{��k(	�!)�?�|�I=I/��e��g�WsQ'�'��@皹%�YU7�ۡ�7󑅺�D��Oq���f_��S�dѫ?����X؇��D1�Au�8���׍�J\=Gy<�$پFHk����S��Z4�)\_X�؅4�G��t��sax9$�oԿУ�:�\?�S��G���a����-*P��X@���ة��t�)�m_������#�6�  �Z�hEx�-q߷W��l�%m��\��-OҬ0g_�I[<N5�f���
z@hŗ��Q�@O�
��p�$�59r����'��m:^kPW�ɦ90 ���	d;}&��)�R���1��E!?X`_8���yL�e4lᆫĞwҘ���y.`�CN�t_1d
�J����
���Y����Q���׾D2����|�ј����W Б��B���:��Z�
7շ�)�b��\����ۂ��80	��خQ6@T/#<���?��I��S�����׹[���h��f�nV�p�o���u�B`�9Xy���&����?0���7��C��K�O��C��O$
o��'˶!�g�T]���B�*��6(�Q�S�O1ݒ�vR�B����r����%7L��mi9�<e�~A�����K+��O-nZ��ou�>ܦ��mv����8ҜkÊ4�5N�-������)yCҾzS�`��hn��+b�[�*�&޾V$d�E�a�?S\h�e�4�'i��}.��|Ƽ��	�&6K)'�pEf*������fM_&�t*���a7��O�a>�R�*�� ���抠�%c.<����x�*���~�#}-PLp5�؃p��5�V_2��٩�����S���I�(��F�$�p�*j񶰛&u�rP�-alwM�r���q���I�sU����s����Zf0�����#�� sj�P/��tMi���b��<��R�6�-^*I.(���ŀ��bv#4���$�;8I�^9��]Lդ+)@�-�����������R���;"�%��t�,�`� x~����R��3*�G��L�u�$��$/���"a���
�0���U�Sr�(�Qh��[	�B��{�~��+X3_E{~Y9�+�^���?ۉ������;�pI�?�c���M.��@���A���[}���*ZǕ��_ܐ#L1��=�2���*��M�F������S,�{����4Q,Vn�1&�S����M�_��1>;)I.h�AL�e��u�L�q����/�s/�
p������&�/�}�����CEV��C��CF=粼��V9�[��(�f���Δ�F��S:�T�O�>ʀr����"�me`��qۥkw����]��f������6�ǒ�*�=W�W\v����;N˽X�!}�s� �xj���.y+5W�92��U�Z��-�Wn�. �V�P�-���(Z'�ˑ&������Q��k�QW���j��	4KL��T�����/���������3)h����+�'��$���.$g�k\�FP��/��2����/Z �4��sQ���:5����䏼��'�'#����P��㷢9p���O�S)��x<|�P8R�QVe�3WL� Nh"���b@N�^�1g�Iȍ���fpaR`Qj�y�gZ�w��(��&=g�.�%���n%���m���3�����U#$��J�}p���]'eQ_c�#�h�Y�2ZH��	^6\A`�if�u�ֶ��=��kDt�J��S;��
�g�� J��[���v�������JP�e"��P�:`��+�PƘ��B�X�3�;F��:��_���& D�d*;�O�'��O�PhrІ�r�]az�v���e��6�T,��������6M|����H.�D�JŦ�ONU+��o����3�>	b�Hg�+�ig�o��x��.���Yk�j���E|u��j�wb�YS�o�+K�h��RL�%�Ps%�)�a��&>JI�'U�[h��.!~a-��g�΅����L�a��v����G���J1�67�����b�5x¬� ��8JB������E_À���
{A4Ȉ�1=�BL�
�]����8;��F��q_��ȦF̂���Ma_F	|�'�n$��(�n��gk�1%8}�/9��&T��`L3�)� <ە���U�B��J����b*'��Ls}1�l�	�� N���F�Τ����H'QM%�\����(��qI�@���ZW]8��4h�����K�o�[�w�k�OVɐ��{�n�~rX����vd�`��;<3��'��8yiy�L��?��ĺj]��hnJM���b}q�Om/ ���2�ϒ��$�M�<� ��o	���Drx��O����Q����ź�ZOZ��
'p�E	{���>c��7�f�(R����ƹ����_�s���0������dܶ'$b����3ۋ3�k���m���/�o�� ��N8�Cϯ��wG���n<��+s0����d{H;s|CL���T\�y����}�z��$CQ ���y&�0�i�35�^�wr��[��3"�PdEsa5�@s
�-)��i�	E�@��_}�A�7�Ĭ��5Z��c΅HAc*>,�*��L�9�*�����&�ֲ�y����N���y�)�q�	�Պ��T�ϟ0$��Ҵ��]�(�V��~rK����ݸ�1e�]�_1E�c-˛�τO��T6�{C\{{���?i�/��"��Zbk9C�W��q�a�F�#q�1���F���d�$X�}��ɹt7}C�$�ڌ���̓��nc��!]T���S�G�b*�~��@��CC�܀,O3?�+8���zXw�.��A�������הJ�������%�B�(P��s9Ո�;:~�;�I�o�ܜ�t��7JXu�:�H�Mq �C�8 �	r���N��˶�,-4�Kc���N}d��jIO+� �B>%;�l�����؞
�P��H6��ٖ����:�tj��qvX��Gw�-���d�j�ZZZ#.iJ�C�P��_5�!T�~����&�(�P �"����UV��A����j�͍�ASo�sx;�
�8���LBI�%��5R�>��Q�8�NJ���X�|�|fs$o!v�F_hzL��آC��^���nT�h+S)�l����xr�cq7l��*��X�g<�$mQ��?xJo��
���8��QQ)�#Kl~ğ��T��������#=��D�����p:���������L�.>u����u*@m��o���yh��co��`�.g�zƇm��[���ځ[�W��A�f�u:p�n�r�D!�$;P6C�y�>��"�b�����skt��@�	9��ꌏ.FuQ�p�Qu�HjQL�A�����;����M�4tE}}QBH�{nh^��}�x����җ�<�7o�ց���f��w��b��_{����D�hW	�<~���L&��8�)��h9ގ�~ �Mdܦ���W4�c��R����~,o���i�1nͬ���۵�{'�k�W��kOj+@���}f�W��se:�U����f�Z*�V�� �K�7TV�r=ǽ�4��.q��a��������<L�����MC5t��=�4�R�<5��?�$�&kE�ޜi*��-P"��ESa��x�&���<����XZn�ƊK���<�$��޼�ڮ�eUfq�j���&��Y� �:7gױ1}!��g�d (��q���'�T{����b�jn��"K3,0a�4�[��L*Af\�{����&�q�m�6��?3���õ��f{�ա����g�cB��B�<�Ӆ�r2g��5^����I2hk�t�T��i�k|��n��$|;���5Su> ���W�BH�k��Ux�o8\��b?#���`�ٔ0<�r��ޒ�{f{Ku�5!&<p"��:Op���|h�P}�Ջ�P���Ɵa�^P���6��r��!��pթ_~�XO��lGL�_]�0A4CA�6���5{�k�^(��ǜR<?�&�M�Α��T��f[$<���c�HC�x����	���e�/g6�n�������
��HSL��ƒ�O�\Ȓ��1�����H�>qɧ�Yk�4�[�R�ܫ�W��{�#l����E���V�����0臙p|�!�G�ui�:,���4����ð��d�4��}=� �$44 	�ӬmL��YD�V��DS|؞�v��@G� ��_Y�F��)Cց��C�
��;�����c7�>[����L1+Y��]�3�&0逐/{�4�he��6�CͿ�l�6i��iG����%����C��g�Y��v�����PR/!4�ü�fy��I��iBΰ��L�0��Қ��%��ҟ��`��it} e��o�� &�a�\�-�$��i5L:g����UIP���f��/�p�n���az#}vb��E?G� !c�l	\���
)q�Y8�\]��(��z�|Ym䇊R�7b��4��������kU�*�i3�?)CR�ڄ<�7"�}'E�㜴1�5OT�|V0���;�R���
�Z����bO�q6ei�\p3��hh���J:��>�8>���5E.ȣ0AS�y����9�a��=X��4醪�"	m{}/��
�{"cŬ��؊C�gn��F?S�lC��.�7������	��*�.$-%�3%���΀���?oo��jchh��9-���|a�`�}�NZ�Ѯ�T	�Csk��q�~�Ԛ�H�lZ=�P'ƞ]<#L��vx_�=�'�;?�SrP*�2cw�"^���W���>k�U,}}�):��S��܏WA�$^p�����̚*�UIq��!T���%7���췙L5����;�Z�JN-G��L+k��lʭ/\`��2��%o�qP�	x�;�X$�ܨZ{���]���#�l^�	�k��a���FM-�.0	:4�̍�wX�_n�E��
5w��7���,/� .�.����W�FaS�b�4�dU]b9M���/k�|����r���p��b���%LVʰI�:���/،�OO}P�e��j��2�>2wr;��b�zJ2ֽHB���GJc�E�⋮/��H\�,�a"����j&��e�1���xH�`��4PD���%66-Dp�tu8ݗ'�)s.�~����8[�n�f�c�7���Ս��A?���{�8G֓�6)v��Bbp�(J	wF�����&���`^4��"~���A�%����5�.w���VJ�A��0��	�^[9��>}����	?p 9��;��Vz�z�3JN��	'��0����E r��0�\��m���B��,NH�}�A;'KS�d̛��͵�e_��,�oJ�G����\�ԫ�+��P�K����gs��4�:S �A������y�A5��q$���B�ü4D�5<����ԎP�w��x�
07��.C�h ��������D�������Z��]�����S�Y���z��f7�I�.��e�Ie���p �ʨ��Z��k5���
Xoq|�j1����J~��	8��r�f�>���Q_�[ɠ�Q̅��R�9�b�^;u��O��|��mut��H�	�<r3��8R��#<�V1c&s�l�Ftr����"]�f�n����̳�sm�
&@x<{*�͠�#�/N:���ת��b�W�迴�:����̼"bӀ�x����#�1q���E)v'���*�4��#J,����˶��f5�j�Y��A�l�M�hͲ3�S�bx���U���I�h�L�0*&(OK���E�J��j?_�xAR��6_�2�9+)���@;��r��a�����X��2���������`�Xj%�;���ѳ�����@s�qKo[~�Hv[h����~�^{���r��*&i6�`{��:��{Z�HI�(^1����g�K^s�k;�h��u�^�_�k>��X�� �~�!ӎ�Aъ�#sQg������O/����fR��md{&6�pDw�z��QA��V)��G洜yk$A?_�wt�7A
�d1	4����c>M���b��f��}N�U�OM����K�UȝC�r���w�LQ5� z.�P����d[d]��R�{��ô��˕
ț�i�����G4�=m�#�.�L�ey�������FpI����Ўe�����W�7|['����j�W���YEf˃Ki���'i^Yn�38_m����ѽK��7K�'6���+���,�/��w��zV'5zV��J+U��|����y\�g?�L;��i0���������Wǋ���g-_��3)�C���}��u��YI�I�oi��g �f(2�z}���նX��aAx)�?٘��؍'�.���ۑ�w�v\v`M��Q��M�P��y�����>pej�Ʈ�8h����^��?�B��N�R��=�Y���ؑlC���;��ڢ���A��X>��KQ;W+���a5��%\6��"C��_`9���M|3������. F=���\�=lu*��"p�qvq����B=�l��	���Q�_c"&�t
s��B��}T��^�t��8��x���_k�8�"d|%I%��k	��M����о�Ap�z����Ih`ެ�|cg���L�����|�'���U�ď.U:K�xE�Ot�xuUs�\�Ųze�&� �Y�}�eW�����`�{>�#_8Oa<|��x��ش-E�K��c��i�I�I|���Q�.���5����xNR)�ۇ������x9����${��\���� �`�	Q�NL+XI�$���=���s5�	vV(Zw΂~��}�훯��,���;��J6ݐ�C2�����+R>��D\zVPv-���a�M���U����r��k�q*�n	Gݑ!(8[�M炪_|�1L�)�#�R�|��lF�������[��79Ha�KI�Z9���;�S���~���u ��W��C�w�O0`,js�}4	1w�	�$u)�.�B��3�*�pɹ�8rK~�ު;��F��y�����ߡ����L�u�"l�fS��\[�<[qg����]�Dߵ��͞x�0$�Ϙ�`S�|/Zȭz�+2��nM��h��`~�,�*�X�뱏�����P���<UZ�����P�/0bު�ڂ*_:�HS�*e�$V!C�ԕ��W�&<z�v�&E��N��cfkq��4��xc�?Y|ݞ0U�Y��	�?AVh��h�3�Ѓa�=�
��J��<Ѹ�o���o�lB�&��HG�2uEe�O�Di
�3iM|�l+?)GP��Bu0 p��8�Z�T������Ԋf�>��\����{���ح�wJ �[\�g"��Gr�u�����Z�� =V�����-?�[��q��wy^W[E���F Z����M���K��'+�}���E��䛶n���s�m[Db�qr�z/�����1�K`�|�/q��r+(�]r�v�}H�Q�sA�=Z �Oߪ��cj��K���z���ɵ~O��mw}x�XK[%<7Ȯd#�D�_3�w�ֻ](�&��ޝ�pk���=����6Tm�ш�ۗ:��=+��^�w[�LA��������,�N)���'��E��Ţ(�)=k�jWi�)4�o�_�Ⅲ����?_[��O{�M�׶��=��LR	����A��#�y����n�,�� 3A,����\h�>5��� +��0o�����cWA�>e����5O����4�������O	�du���ao�������7��5��}+�%�A.�x5s� ����_��	G�h:7M�&��i�59��p�jqq�O�ۼ@�T+`E���w�?ow��.��M����[��3X��8��_q��h7}����b>8|�^�=_��
��H�i6=�z�C�2uCa�T�����(���(�aM���4ѯU˺�� M%�ˤ�c���V��ތJ��%��ɐ9����b��zg��o*�6�AK+��FK�6u�"� �k&�4$��\(Y.�Mi�S���P@ȶ�$��ۃ�D�S2�"i�?���nl^i��U�/��0����c_�k�&9�����*��=֓Nk����.eyx�����=��LvK��Q "�Y�x��R����t�B�[i�)$T�[PxGv�V�Z��|�%e��)6��՟�G`'����edz����wn�lG�����ϰzp��Ǭj��2"b�*�R�N�/tG�(�,�~�5J7�u�_��z?]_�|@��l@�5M��7A�M �W�h;�;eQ�:�b]%�m �r0����D'�����.r�'+�k~�Y�XA��&���^9/.,�	��C�z�T,�]��q<J'��ҝ� � �����o����k���Uy��u�>�o��3[�z�����ڒ�XBuV�mi�>��t�ymRٟ����s��o]ͨV&�	�_x�b6���j��V��hm���αr%�?�_��N�����T���UMǳy��[Y��~h�O � �E��M3�B�_ƣ�kR��˶%��o#��9��5�V�D�*��e~`�FI	�3��V��kJq쥺��G��r�v�f���'bR��H`:go�<)Ã�5��\�M�N	��,C���7�)P����pC��>*��CS��S�:�F���_�Q��{]��ӂ�y�L�:�x�K�������tJ�vX��:M��?9�r�����	uCe������tS�f�r{��`R p}�̍ �Q�b*�Qna��ޣY�A�q�#2k=�������l+y��U t�[%�����J����ӂ�
`����$�1lP�g^q��u}^Cl�;��VɆ��:�%P� }�hJ3�?8	9C�gs�/9���4@�o��\q��N`3��o�H])����Z���+d�bꭲ�ЊMMe�o��e\�T�:��C�j���G��"�*yϙ%�*F�@ʻ�ҍ��&�Sj�G(�tl.�˕pݲ�u���X�2dHn�p��9?l��D���I��A]S��[6��o��N��Ҵ@|}eB���8r�w�ʾ�5XG�x��d髎�h9j�xB ˥o@���Z!0��E�Υ_�׶�=��2��3Ca �мS����,�2�D|���Ou�"j'>ZYTd��rY"�qi:9��ß�5Ξ�u!��(�f��[c* ��%=o;)�@m�����[��׷�9�1$��H.
��x�/�& ����g֦u�v�_(ak��%�&��DT]d�Ѷ�[�cq{ި�oo=�.��р~�-����ѿhU�K�ժ�ie=����t}�AF��vqZ`�6f�e��{��(7�jF��Ic��Z��&س��g�m�!�4��S�N��R`��^-�1��85�.ʟ�S�G��"�/r*�g�A��כ|k�E.�;�8`IvL�����qu=�\�"��B\��d�@��*M�1̧	�����3Ŧ�UɡP82#�l�G��6����V�C:��e�*o�s���\ة����6H׋-٧ݗB��IT�T����@.^���q���D*�3��D;��3
"�W���(���F�|�;xe�>VgQ��cͣ�1@��wÂ�Q{֠�t�<!�)�_�����?��Ŭ��y8�ٺ��WMǿ|8>���4%V��+��xT�9�˴��y)t�����"!�\��|XX��д����i��y���{�i�BAC��/DŌb�mK1�� *�Ԕ�	�,� �&&���t$�Õq�xr+��]�,�I�H��������̟��(�A���bt/�p��$i�N��F_��&�4�R��V_�Ƚ� 7���X�Q�wk������ϯ�I�0�8]��>@��[���Hu\ ��W��8CT��M)i(����P X7{k���\������n筢Ʒ����̪����{�1�^L�9��ha%I��K�O�OɅ�Ʊ��=�W7�l�I��O`�շ"�l]�yN�-�:���bH��ߦ�Z숦�E�����|sI��>2M/�&�M{�4~i���_*�0犙��,圦rwt*\���R�<P��_�ъ#6J��CNߞ���=7s�����P�x�ĕ㓵�1�_r���D��
zҨI-dopu1K�%�5*4�򏊇�qCe����}�?j���y��C�Nԫ�������_���8Ԟn�rK�VLͲ4Q�f�w1���l�r����&!�����ds[L�h�jGn-�Oo�?��S_"a���VgtDߒ��ܭdtK�Zy3�w�x�͵�f�X�������y 9��J��HX1=u��[�x˃ ��r����'\�,�����;�I�y%B�(sO�n{���lp������ ~B+���Mav���G�:�p{T2��\���c%=4��C,z8E1Cp��N�k�5O��-���|-#Υ�?�+�^Y�c�=
�57q%S��h��]Q�W���V|�����f���.�K� �hK2[z�/vOyo�2���ye��ɶ[4�)U��]g{w���nO< ��K&&y��i�����䬰)��e,9X�;�\�m׿�>Ul�Q��"�{6|ڨ�>&A˝���n���u�P�'O�h���]���q���_NzW�8���j�[��|빏��AT�u��Ԃg[��/T��u/nJ	���*.Q5�&g )�8�F�ڗ�!b�:w�h.٧��+d��8�#+���}5QV9Q�7�PW@�W�L���00���m�G	�x�lA����,n�{�{͑�)�¤���o�-{,?as��;��b��n��7�R�q�
jxJma�ϴJ>�绻?��P�`H��r�CW�!@�;
��;�͘X�Q�	*�t_�"��{=�����P�A�s�/�[Q��e��2���+�������a�G͂��xVT�d������1�`�a/�w2��o�HAl�rqd�67�ᒿ��A�l��U;�3|��O�̈"F���	-�UmLv�+��,�`h:O���|"{�ON��5Ub����خd�?��;jگ��.�U.�qʍ"0�Z'����/��ۺ<G��z��vX�@��KWV,�~a��q��Cu��T��J�od�C��8�������0S���Cj�H�Ar�܈(BX����&W
����e4����x��!N�[/A�6t{�l4��6�B�j��]ʱ�[E|+YH���E����m4�+��$J%۩E(�7�
�����u���.��� ��T������ٙ��eE�<���w:EZ��ږ�q�*���5����:uP{�0�6���	�]���&���g Cf�y�e� ��cA���֦��v	|L埉`� �G���U�{R~�Ln>Im� >jp@�H��x�m���p���|S���Cw��PP��f:�ܸvw��,n�t��OBaˀHr���z<�T�2h�+:�b����e\�V��+L�-�n�i��zH3 ����y�MY�1G��+y������@b����ax����޳Դ��3q5��p�=�x��x�_l\��d&�~���lr�^>$ʩy�AގJ[{M}\!|�>Q��K�Fe��sT��N��V���]/��(r;1qƴ퓗U�����>��My^U�U�E�Kщ?W'����Do	�p���o�LB�¿��4�w�������8�O]&X0����xU��-��~͛E����(�p�� ���R���M�~#�-Q䯴�V��;�=�f����s��D��eG*?g�5a�^�RW_�8�&�P�/D��6���w��:l|[֪�ګ���
�t�V�1e2�5���F<�T5m��N�𦾉}���Ha��9�������B�7�1k�og4v�K=E9����4<U�lp�y�᷉8
�/�hɂ�.k��Vp#����ɸ����y��)X�N�w%����h������ǟ�ö��|���aosp,#����ǁ�f��f�6�D~�(���#���z�h�8qP�I
�:F�����&i(t��5_��r�}:o�Z6TB�^I�  ��s�E�[����R��C���B�-`�f�\�ϩE(���9����+�*�;;pQ���ip~]��q���Q�Xs��)q&���v2������@��n�yY��)�GJ���j ��~bn|�p�,^n3�>�EK��7�&b���bț���D2ry��S=X:uٓ�n���'H���1��K�z�0�m$�:G��TF�e����UG�a;�c�j�T-����}�r)A�$�x��1N&8�cz�{�PZ.��[��K)Clk�`���F2�4B�5zn�"�0���gM�'b�5�|Y��z�`�	�Y`���ROyo��r��<���䤲E2`�i�LU�)[U�ڑ�PQ�쏪��o
\2zoH\�BѱL���U_�׎ޞ�m���Sh�0ɼ	��1x$�cá���Y0����#x�������<�A�]mcy���X��]���Zu[��/�໷���/�J+�S��G���;
���`=�#����=Q��{-���B~�-
"l��w��g��F�������B�������Rr��N��u�C?������K��1�i��-�t)���"������ҨnhT�j�����R/���C�9��|�G|����ߍ�t��fP�Yf�]O�y��K\ؙ�
��[���������C�N�YB-h��z��!�Wj������Eǂ��;cIDz�HWg� ����҈�n@[Ռ�%���ܜLϋe?X�s�G�Y��=dVd��_kQ��Zc��}Sw~�u�Ɗ��A�L�K�q_���Ӷ w��0�NL�#R�4�n�j���Bs�K+5�Ɨ����6�H�k5�Q��E#1�c� ?mz��L�8���5=��"��IqHQ��u�sc{�����D�6�E=R[ޏ�su֊����NrN�V�u��}�w����D>V�G[���z��1,�(�}�)��s�,���8@&2_%�ya:l"*��y���Mp,��hs�����Br���r�Z�~�wO�V���*��z����E�3o���eB2�)������a"���I�!F�:�l����O�t��q�����,#�U���"a\�uj�ݫf ���_��a>�ߗ�����[@�w;:0Ld��ӗե�yrٖ[���*t�>ɩJ_�)e�6.@��%oȼ��|���3V�B�}�W~���CΨ��x+��z1_7��`���]\i��7૫�����V��)&��v��g����!�����O�o"�-�nU�M��_�4���s�C#
��g]I��4<�w�"�����+gDQ��3��Ī�&����( �s�%�e�k��wd����H�r�}�}\[t��N��J)8T�;i�VJ5%4K;_�A�+�clĿh��W���ڷ6-�g�J�[X;�8,%;wO�@ b��~C5�zzu�/�[8+fc0M��6
 ��_j35�=��$�p���<��U ���7e�|��S����,��nIP����H��N�`�S��3���wg��\oZ�g���i�L�eI���G��9*��t(p�����Nt��Z^���$����� �-U�����y��k�)������s�n�ω@%�w�S6�@:x�gǵ7r�N!hk�\���7Q�)}�kw�4>�%��C�hF��d.�@*�|��vl��;���w�b��O�,�Ӎ��99�{⩜�YJ��nn���:O���g�g�u�'�x��v9W��k(����nsGaO�gb�x�v�6� J���O� IJ\�%[m�ѳ�t�U�ZMy>��8�K��#c(q>�:9�����po�O6�[���l��Iē��UFQ��;��g?i��d�_�2a�zu����mm�F �r#�!����&r���(���Y'ӝؠ��\ևq���3�K��,�����s�5��,��T7�>y�uX�X�}Cf?�����}M�\[_�'N��
�7�v� �E=�'m��H$\߭�i�G��"	!��i'�L�o��@��Ü�!��v��G�A���X#S���"Ҡ1`�-K*����c���J�eV�L�0$� �����m���E��<� ���c��q/���r�$q_�u}b��_�ߍ�UOp��'����F�c�_�A
,����m;%,CUBQ�y�\�����O��|�	�J��>�m��s=B��A��q��'6g����L�B������2�)08U�T�`������b*k)�P�&�t �+�\�E� +���m�-5��{廦r�.Ugp{seS*��ɘD
���V��kɜ�c?G��=��4\���G؍�Ox�)��!&�i��i�%��V��Z���\V�U9h&���V{�(�*"�R�Sc(o[R�4t����lqC��,�银��&��A;W��V�.�����`g�W���m�H3ˡ1X�m%x��l�6�2	;��Q�`��2�;�e����׽7����t�L��=kE��si^��َ�	�4��#����Me��-å�p��&�*��d�ʘ&]�Qb�2kR)J�U{�P���@+�UH�b�z��@K����B�P�L�Q��G[���'��dě�YD�˅IF��au8(������_�)u�ݺj�r�?(��j�W[�����çz�]�Y��z ���],���xR�> w*���V�zUg�](j޹�YL�p��㏺�j�<����$a&�yn-��;���˂���p9~�f�p7Y�}Bz����Z�2<ua�OX��}��50��s!Bэ�M�.�G���1�]׈�NU7�h|���-�.kU����0:
~d�rY~w��4AX�PP��5�͐��8��^�W��*����el�MeN���d<2S���m�@�;��#0x.�f�d��@��L5\��h���I��t�2��t2���h�D�g�A�-gvq�#H�d�9���;�Y!��W�P��j��X�f	�:Q�-��yj*Kr���+D�rߍq��Wum��iPТ9e: ��B״_��bQ�Z�.��"�_�1R1���	3������'���ޟ~;7��l-An���cK��-�Z�����զ��J���$�E��ĭ���_�M�9�ڱ ��A�h_B[�r�ůɵ��h�u�=vL6А�tAdo-�P� #�׬T�\��z��bA�`'��xOJ�P�<_�!롯z�������4�:5;
E�u'l��E��0�"� M��.z�>2�����
�h!z���qi��6���-< ��I�w�;a�`�=Y'��2*�a�ES�%j�(��sb)�<�+���~jgi�7���|~o��{$�µ�d�{����i�� �2@�)o�����tC/�[�5D��_�K_�/��޾��<'���v���|��`�S%8��!J%3]�I�}Cvw� ��A�X�!���Kۘ�4rܐ��E����\����(��}WZ�� =�P�̯R|��3�JF}t<��y�s�/�sD��Q���SkW�&�gv� ���iݴZ����0�SԍTt�g�m����_���.JM��CY0I�s	+(��Y���~�0g6�,��2*{��,�d�;\I�+ݳGQ�A����h�=�����\�p� �~r"�jWjm~3K#,��	ۣ�Ęq^4��k�6U�Ts�
�3;V���.�R^�r��{:�\wV�=�w+M!�呆V9Bl��g� !i`�?�����P�)¡%Q���*|�@�Gm �2�EڭÛ(uA�����,�-ۿ�yR�3�*�5W�z�4Fds[�ڥ񶀓�e�m)���:G�W���`��x�O�B�H6�,¼��h�^�=i��r��&R��W���=�)�:|���G�!ήt��:���=�v�˕��N�t�S^Zf����0�X3m�s����a�O��U�'-��A�e�5\�Prr��|+����'���Λh^��ŭLcO��<2L���F�J�Ä��|��eQ�ZnNC�$�H����E����m���������?�t�YT�e�8O������"PP'e�����|����ܚ4�G���۶"&\�С����aV�%�Q62-�j<�)��4T�ּ��T�9�x���-\\�a32�$�sb�#������˪���d����,"J\8�^�.߳��$�D��|�T�	Ѵ���]��yIK@�\W�_ڴ9���i��j;	הm�

�m��f��"���5юJz�su���z_�1��3#�izy�1���}��ZJ��~�Z�?*���Qų�&�z"_C,���������TO[]�C2^�r[����^��t�x7�; ����n�h�V�'q�kV�z�1ڐ��׎:|���Z)!��xM�P����@����D�v��@
j{
����r�:f[�*C]��{p;�� �ՇE8���+���NM2kfF�]�oWɖa�I��+.��ȧ�ާ�^�ghc����H:��ð�%�㞋e���=O�����˚Y�:K�.���{�8���v.�@�������ڏ�L,�"сvnqP\�&bğ�0�6~:�Y\WM([}���6ĺI�Y�[��n<�b7�,`J�ג����X������ʈ�ϳ�*�@cd���۔����\��6$�D��Y�c�KAN���k=�D'�#{�z<���_����sb�"xB�����N�i��4WR88td���2@��2�~��]���ю��u�l����J'�}!�F�2d{$���p�Mj��3�1��g���;
j[}_Y�̵�ų�,3bN�vþޫ���%T��鴲�kS���h�H!�=8l?��Ll�i >{��'��~<��H�J�ˢ�'u�ԃ��c�V��NX����w`�h��mg�J���kض�p�)��J��l�L>�����,��� �	��#,0�s��MA2�u5��(�:��o�=��,g�U�I��\e���G�y2�}�hܩ��K�E���YI�M)�r�����E`�	ة�l,v���A݁�6\�m�_�r;�jq���]t���-2�Řప�^��ɢ����:Է�LN˼�>�v�+,&�$C��=ԉ��G)�pQ+O*~> }Ww��L�$)�P��r�?/�_������P��8f�>�l�L� M��7'�v1��+��?[�UU��Z&	�j�B�s�%��wCxo��0-3��������^m?O۽��w�\�wL`�f����>�j4'k�@��C%*� �|���G���J�hObZoZ���U�j
�+�B�ePq8U��~��n;���Wsu��Z�頪^*g�k+¸<{�]�X�
DWs�a1`>�J��׍��@����#���^�pIGA1Q>U�	Hj��/U�j4�;�r))���d"b�b��҈WҤ�y�ft���krFs�����k���Z��v�'�ސ�  ����)��>۩�.���=�PUH������,M@��pn��s尐-�Q@�֔3y����ntv��sC�}⎞<a�X�#���Q���~=p�E�p0���5	J�
�����9"Q-�Y�ܝt�UN�z��*yl���Q��T�@p]=��Z����[����u�;��k7���m���6dkY_հ�&ʺ��sM����b�j׆�W�\vI�c� Z�↺k����s�A�g�{���)�Z����^��C���<!�}�pUǤ�̉Q�|?1N�RbL�'�q\�M��T�]%f���9��Oe�йU#C
�,�����ܭ� ͔_0q���[*T�tҤS&�[�������f�S� ��.	�nɒ&����5�����X7�7vK�4Z:�1��	%�{=�Ɏ�5t��~7u^B�Įض�k�\;~'�d��Ï�R>YD�����!r}b�����]����蕧F�C���ӷ7���Ƕ�5T�Ez�{rw��y��ݪ�x�:��m| $�(v��־�T�Xz��~�孙��ܙ��CNũJ��ڎX��ǒ����F�̩�#Vhؼ�QV�uF����Fu�4q���?Uu9�[q��?��YX�qC��W��é���LG���tDnz%s�|��}���i)l�����6u��+N�~\�n}���F�:W�\�0y��l���~0Y�<"�t.ʛ;�}�v�
��@풒�o�	BbZ���'�z,I��I�q P�ç.�ņ�;�c�z���V��~� k�c�A!7�"�C�E ����w��4�i���{g��e
�sm|LR2��q�Q;ӆ�]b�Kͪ�Q�����������m�����ۧå�-#���6Mai��ux�$�A�XG���(O��u;�"
5k�����P�4��6��*�eN�iq��	��v'���r�5]P�gc.0�DC:���^���{�A�7۔t�OR�3�M����-�9Y)#6���[��&�Q�ܫ��:�6gg ���k�7Q���E�mx����U�ⱃF�TiB����#��!��$G·��-�k���W�R�*�N�Di����З��DQ��xC�c:����Ƃ�էK|��p<�;)֚����t�����^�l���L�* �5	:��?�/�J�������y�ۮ��M���퇗�R�*g��ܛ���f���E����=&�i��|ؙ����{Wo�el�IJ�<�͏،�
��7�	 u�\]���nm���m���ԍP�p��#Fx�[ǂP����'��y�0؂��� z8V�*e<)��_8-�b��C�n&r�;aX[��Z�{�[��2ܺ���Λ�kq/wR�^DA�1)�K�q]�q6���k��$r�/��и��aگ���@D2D�0x=B�TLI���=!�ö���ԡ*���D����Պ�|� I@�SJ�� T/1�g�Y� Pӈ���*�4�oN�^]�y�IB�>����Pw����t�Ϛ,dI������EWN��4�g�mc�Q�.X���?X�-=v̤��O�C+���o��X�W4`��U�9��I��m�����qQ!X�s��V����SC���5D� ��3��I~ު���l޾��hmϳri�j�@%��8�%�+g��@)��,��[t�6��{x~����bz��f�u��JDD-���]��q鑐��یŹ%��PC ��tR���0J�n�C��ǎ/ڼ��{|��	ȝ64H)��y�,svܴV��g�t{��0��=Ꙝ��P	�K��b��-�L��:��lY	W� ���0ߨ�_�ɋ�a4.�M%����s_TԒ��g۲2�:A�B^���V{5S ��Z��]�J!B��j��|1�cap-�$�7���E���նK1�q/�J	�F���=5�:eӷ�M��<Ď~���ri�
1)�u��Np�ң^���iǩ5��ۄ��=�?8YUw�\ů:r-
�����m�7���`	#�MV��}t�0���FAL���g��ɏf]
�wn{�{��?
���E��-'�e��c���P#
�
�~�KT���y9d�Uy�	��;��\����:�\�1����1v�����ŦI���3���c�q39�3�j~���upI8�wxF�����%5�>�ӥrv��u�Z��B�əq]�{���7`˶q�� � 2"���{2�ꥬ��c-}���f]s�7-�?��\����"&�:-K��H1,���ki�K� cx���E��)�-[�ڵ��.��y4�R2�A�=�٢�+���LJ�����lK��nI���X�(=���!�~G�<��A��YTws�%�i��,Kf����W_"ڱ�oכH���T�60�֤ڇJ��&���	nw�>�ζ�͵b Q��r!'��/���������a�<*G�1�ӭ$�I�V!�wJ/�+q_H�o����#t��ư�-E`*�˘����$	�ͦ>�"fΔ�Zu�U��Y��$��
��٩��f]Z����k����>�[��T�M���W���-М��'ڔf��������׆�X¢��֘��yrOb�V\Y�!=4`��w����M�w�w��[�m�5?|�_~�q�S氄��F������y�YƢ ��üª��N�Y	�,�BEj�	��P��|��^�:~�1���jE�.i�d��P{�~櫣��X��э�e{"@�2i8�a\-�zR�꾎a�z��ֽ�1}�}��M�t/)�b?���{=˸�N�O}������?y���a4�~|:+��K<��~u(����pV�M�6M+$�7ݟ�38���B��Pn��p,疢�_��"գ��+�ϣr.b��{��F%&�t���nx1pmW�0j,�)�BuS�{�������^P�>�?c���~|�G,x5�u��)]�x��wO����:.���Sޜ�AFg�0��h����<�>�����n9��q��~��u���Z���槲�dp�U�o��ٳ��Q�A��ǁ.�*��N��aN���Uy�W.GlÞ�e�U�P�-�3��' �Q"��;&Al]3t�N����NUFz>��*�N�;�m!�8j��;z�v�L|{^X��yL��v���鮓�`���_�'Ú�����z��>���	���w���<����?�hj,;5<�A�����|��B��p�(	cGT�2�A�!���E�٠yV�ׂZrz1� �S�`5�Z@[��22Uʹ��{��!s��2�5����o�8*����^D�8�����8���,�vOn:��fޖ}�J17}��J��	�Z��G�"`��cXgw�� ��9����B���O(�B]��R�l���Jx�]B�����~�^́k��4�4�։��:R�L#����V�������>�o�,��/���7O���Vp��c���]R�r(��|���o��7H2��b�`�[��ߦb�e�*ͯ	k��z�����|�Z�8��C�2��DOy����O�V[���!�Ȃz,�[��?a�-�sil�h�O��!+ Q�?ɣY�6aes��@���������|(���W��q �ˇR�[�Lu±��ӍCVYx�bPĜ%�2�ڹn�ܹ�v�K?>Wư���2u�{2p�	�u/����"j��Bk��J���`>J�U��;��:$���pe�����=�$��bxT.���BG;�1{&?�5�U��,�c.w���K��ӣpz������a�2�ss�nȐ�M���� ��	%�{�0S�r��rY��Yj5���zY�Q�*� 2�pN<`�
'd��$,=[s�(�ܰW-.H�-i�Uɴ�@�%I3�#ԗ���yD�ѵ> )�L�C_TD*Tt�@0��h�唺�T&F���L)��"[�117�X 5C�ӐZ7h���e�0��l ��ǝ�Za0Z�`rR6�*Φoo���<2R�#}z�\�s܅�c;�/��B�Ol��E���a�kd�T|i蘱�����tJ�k�d�R��4�6�����A.;��Eu&uH70q,�-bZ<�bL��1n���S�9�N��X�N��*:� Ʌ��XI	<�͉�WLyc�y�D^�E���,Q�(��b����3�GF��ޜ�=��O��0�)IKi��=[�i_��w �4���9mt�pI ��1E�"�j\%#����/$���Μi]Nv�"�E�3����&u ���څ�yøe$�cn�����kd�3̫^�R����?���_��d���-�q�!c6��bw�*�beCQ��+�AV6_�v�+�1�:�]A�U�ݍ<�V��5]��m;[�f���-O��|��`���V��S�L���X]2U ��Jȶ5��Ѵ/ gs��Z��6�K��k�U�P�\ƾ��ߎ�{X��1-�c�m��'�BqY�gq#�x��Q2��b	`TG}�°Y�EV�9Qg$���_B�Ů���j���o�ɻ7^�9�Xw�3�K��B�mv��R��	ZLY����!��{A�\�˖������<�l%��yq=j�fQG�ú����zZb�f��_�7����1A�`�*ϓ�,.��hcZ�V�����>*|�g������;�R0��ڝ�@���Zg� �|AQ��{���5Z��zv�e�ՠ�����J}��+ǉ�D�#�c�^+��td�<�.���L�0&X뷝����k���	9�R�;�X3$���@��{|�O�����a����W>T����:n-r ���0��r�:-�OZ,�1Z������O~�Nc̖8S�	��2MM�3Ko� �,N�?$���}*.`\:�r� ���Ձ�{H�Ae4>#�A��kQ2�ģ��ӦT�(�a��^VA�+Br�0�,i�F5I���j�?�'�prᵚ34Ȯ�"�_��<F^�O� ��b�_�wKR��[;],g��]�r��+@jM�Y����ĠMo}���m��� �g0���� _ܭ�X;N^{:��Fr�Kc��Z�tp������(���g4�q
ˍ9��=���<��
˒�r����K�#�%�U7�Os����1{@.'�\�QgK�D�s�Y�5�^������-N#
7cm�q�W��*wםB�FJD�� ��9XzP�츌Eh�Ǐ߭\K�s�5/�o3����E�<0�ܹ�����n�%4U���d���c3M�lXi�9v�V�n�\2/�Q#_N�&�~�AG�H�0��撇%͊�h�Ӝ�j���P�7��ϖ�M����v�c׼���BB-�g�>���z�0k�?���#�����*_Kɑ��]���b��a��P�`�7S�8��
�)˛���<_��}�Ы����4J�T�ܗ9�`�Q0.Ş����1���v��K*
:.f���J^�P�ݯ1|N;��~��n�aE��t�-F5�}�އ�'�3���Me0<��^�,��k�	��9�IC�|�O�Uo�oSc�zK)G� �bR�������&-��lHS�X��ڌ����������-I+��|eV{Uh��
w�?�ہ8�c^��^F��h��MJ��K�Ü$*bv��R����V|vqub-�[�D,g���|��5^#�<RÞg�
��1v�X����T`'|L��6@v���OOcì۸`3����y�X���J-u���m���U�*�d��P�GH2į�G�cʗ��?�V�N�i{yt�k�H�,o�~&R_�ƛ��2V�r�*��c0�P��DN�����_��U�h��{����rHg��m��Wq%�����>�?��@d}r�]ê�x��7�[I~xB�`�����6$5�N�ڗ��bz�_������:������Z���CW������
�=S��auy[�K�d>�ORr�R�q�w	i��F;�]�3Y��Zy&dVg��&��#K�%�k��V���D��O'�q��A}�{\x�7��տf��3?#ŋ5�����s9<�sP��)�������S,��6���<�"�낳e�n�}��>{kD+~u'r�ֲ`p�g)��J��k3�����^�*�G�|i���( 9�BZ{�`x�y��\ݣ���"@R�A�S�u�p^'H ¶iW�6���b@[��.�Z�o��ZS\`M�1s��թ�zA��l������f�٣���v�u����s�`�Fy �͘�����Ps8��������,n����Nҳ����1�D�T ��N���邱$K�\ ʄ^��r�K�A|Z*��r ���t�a�~�2�a�=���x����#�Ÿ��eWk���y���<U��Y�{E�^�h��*ĊJdd4�!:n�ϗ��f��;�Ӫ�D�'P.x;�C���8��G^T��
�z���"D_�rI>]c�N�s��B����<Bʧ餤C�ǫl�.���1�f�a���2�4��Z�옂������c2i�i�(t�-G���N]=�qh�W�,�`,���ӑ�Y��,���Y	K|}pe�S�p)K��7��뤽��xviA�-m����e����/mRh���G�0���/�[Q�Ʈ�E���"Z͏:k�]%:ƨ�
F�guf=�	�I�J �Y��)��O��Cr÷���U �9U�u��$��?7�n2h�;Mf>�X�Q�߳�THJ��SF�%HL�ڗ�啧��O��9}�����ވt���S�8�H��|�X��Xw��<�XJo_�B�UFBfY�F/����������ǕP���j
,�Q�"��<Q�:B�z�#k����/j�����������J�R�|_@WT�?m�we�M<���<�xJ:
��_ ꭂ9�tc'}�h�r ���|R[$]�;E遀��D�~Zz��m!�Z���b��o�/Ŧ��活��
����tQ#�d��໅�v�壃e�:@������y�CAq�!�66��.y���&D>O��9?�0?��[nT�<e��D�Z^�xǴSX��m蔝�
U��K�{��^͘PXQ���E�C����^̝�σ��d�X�a�S�����$�7}gjS��	���c�N��Stc�Z'��F��+u�Ws��]-�Ɛ�r��>)LC��L���>I �#3� F�ɗ%L�91ź�5 ����#q���%N���R�F�Д�v��:G�#�c_&��٪�5��o���龃��9�QV�O�1�z���2�|u���϶�j��'��?�{I��&K�1�8��P�A�E�T�97��:T>o���2?s��7a����`׵���[�����	�
�{�ܪ�� !�GW"�z�N���łH����Q���ԆR���ē��1����&�;�d�lPb2�� 5�.��s�E�-�`�g�$���׷;�̓=����6	�7������Z
y���h8Y�㧳�ټ(�ڼ�|T����]�0��$ƽ�h?F�!� �aV^���WNM3�;��Ͽ6��O)[��߻����\\U��n ���K�1Kl�Ǿf��8f��Z&�uVA��9D:�i�d�!������F#.ˤI_��,"B������`��x��"�Ppy=Q�����_,�L�����As���Gb_`ze�����%I��w=���6$f����8 ʬ鹛�W�k�����S����9�$Y{�
+�fR�n�I��H�V4Ot,�c�\v`�W���!|h�����/$�uע/ˠ���a���z3�a�-�,h�D�J}��r��4{�zD4���j�}��-id�M�kT΀<�q��y�� f��Bٕ�ȕ��>2MYYa�n=e�<���l�������)'ަCh,��d��R����d9�1��
�SD�i�	OL�Z�9)�As���q[:��IHs���8����s?S,�=Q����H���w���B����*jFZ�+�HN�v�Y���C����F:�,4F�lʍ%$������7��^�v��%Z�J�l����I��`n�p��
�a�S�f��v��u՘8ExY�6:Z��7Q��,�~;Tv�k�,3g;�o<jP�K�Q�$n^v~j(��^|��7��>��8lk��@��b��&Uu(64�&<jY{��7<�1�>�""9�J �p$O�\c �ū��Y�tl���n���Y�6q���Һ�I�΂���xÐ^{z��Jx�I�_��!��R�L��7 �r[���NKPݣ��N�>�U��q6�w�I۶3S>�R����ޣ^CC>d^�C��QZ�k_�����NW��׫����T�m����$�pp��}J9���s���2�� ��e�˯8d�F8��n������kK=��~��5R���7_@�'�> �&���bܛ4`�ud��������G(T��;��&�^�(�Q�=ֲ��H�1�՟|ꁧ��0��ye�'�ߐ�}���.j��!׿���ى��x�dmp����.[�!���A��q��0��=�~&mX
�D)$m2!��u�����Z�#�"�W ���ɤh��uk�-��[���F6��%gK��46�, �홨/���w��7
0x�Wq���n��>@��n�Yj��4��\�@65r@��g���!%{�6��
H�Q�]�1d�|}2J��T��P�� �=���ֺ���2����N�^��DR�#���w�?�8���%���_�~Nc ۥ�.��xQP:i�<|��x�
�I-����f�";�B�Q�:�8���(�y�u�]���s��JaM5z�d^p�j2-$ν�m)��F���t�������^�ѷT��J��@J���c�昬	�x���t���+rvGW�7�T�H+����*�������4�׎��ܭ��MUM*�������sm��Ѿfo	���o	E�~"�A͠7�1��_\K�ߦ�R~ܕޑ���#��_] ��(��D��X��u�,�|����꨽5��rt���MJ��B�b�g�$�kb� T��ĠfiѬh(y����ٰ�_��_�!PZ5��5U��-w�*�Nӝ]�frhy�?/�~��g5�lq���5�2:j[z����3�����~2!�bVz|餪�]��3,��E6����bɘ_K8����lk�����'���	��y��#��#�b�@�.��2J
�kO,Yv �~�"n�񢠞�Z���+�	U��}�����0��%w��Ӷu���s�C�!cgGI;�L�RG$9,,�l���]�0���D`�(g�8;��όC���|�n���0(i $�1mB@p�  h��l�����O�S���7O�(s�^� �$
J0d��c����� @���]�aс�1�3��f�W�^��'�@}qܕ�b(�;����2��,�$�Sv�o��r�~�?r���4;A�����V�-|���s�1��s�%��XZ�C#茜�qrb9����g����	���')`t\���G�6ȑ	����ζb�]�\�7�$Ҹ�Iy��u7���.uKV���9<E�[������Vڼ��9|��*"������h֝�^(ܰE�raEc@���g��/�;�t^NY�ؖ#�bX�g�qX����h�(������x�p_]*�W9��23+_���>ƞ��7'�k����{Y�k(4��rF�;|y�u�=�W:��Q���0V�U�~]׮#e7���{oJ�������
� ��$f�|�v��s��)RH9�����-�_D�ϊ+��݇�|�u��R�Ё�br�p$4K�۱�;������YPO�.���S���
v\���p����m5�Ko��:�����ν0�1
��[�D��I�3bW^�捙f�ݚ�:B���,����X��\W���G<j�PI��yD.�м�g����������S�:f˭��t%��|7+��0ejl=�7�D_U���c?����g�� ��W^���.GZs���U|�e��o���ʡGŚ^�;��ƅ�i�^�kj���$�>7{1D�[�KU�������п�́�F�������G�K�Ah%S3��Z��J���8�G�r�̼�R�\r���n$L��h co���ڮ�<Å蝅<[]*�:��ҁP��ؼ\�'�Q��Ȋg1�$ ��:=�#|%��b��#�ϙr��Y2��~#�Cg-q��]>;TY)����H[��r�vuC9-O�$%S�e��R\(�^�4�Ʈ��!$��߿��)M:
��v���g�o_��9���¯l+kLָ�:��wN+� f�q�O�4�$�VgЈ </���ikUy2�x-V�3��̷t5'��:�lq�Lm�Oũ�8�c�x-��yn��V��
D�\���}��f5�0sD�8��T�_SpH���\��L��� +�8 =�o%ҩ��\M�ey�-&(c$�!r(���	�;�E�MIݲ�UAt��ɋm����}P�������e�
{u�,[14�u����L�<���ag��	w��ԧ��K��>ͤ��U'CiH���@�ᇔ�?�Q(�*e�`��R8j���d^+2�@	i`��"ɩ�p������d��-F��Ez~�	�e�:$��FM�j�k��wV����{����f�X,Ԓ�E5���|ϫ���ϸ2_��"��VI��ռz+�T!{�.���b�p���7|H?a��hrb����{���xn:��P"'�o�d=�Pw��c�L������y�I��g���*�����3��˅e,u*y���eK�7�q�_q��B{/��؀AR_�]��p&OGo�]u�Pj#��~ҡ=F:�oz�S�[��;Ҏk�He������r�Գde��XB�U�U7��z�F�`���a�����]���M�E"�F�i�d1��}XȨ�@�@óy4e��ɇ5�T��.@�꒒�o���A��7��$/��A���v��K�{g;���r啎2[�&H=?�"��a3H�bx��	�_l��S��/q2�/0u(�u�)c�wj�x@_Z�	���:�.�$��!������'���6̓$�y+!7$8M�CۙJ�ByD�ܣ��u��@�%:�J���<܍,���
�*{��R�!1`�R���t6ܟ
j�$0>���Ѹ<:g�c�ֻ�0�P���F�ZW�C� _�"�E����� CS3�_��U��mu~`�XU2f�՛�6v�o%��~o�]��f�~*�mu�#��r�X��^JSq�e�}U�)Y vP�ה�і���s�&-!���/����
�䇆�Nc/�~��V�/����^�>Ae��M;�����"u���@!�NT\�i����F0��֬X[l�{���5�$!��3��k	}��W\\�"f�ڂ���u��:�8TJ$�d��&���f,6L�eO��)v��@�T[� �>s
��O�N����Jʎ��Td��V���������0qĹ@Cg���E}���V�N[�jf�Q��֏U�l<p������Ѳs�#y�=:��K�w,K:/� ��p,L4�t�ձ=4�"��YS��=5r�_EG,m��~���to�d�_],���01X�(�!�:�>.�u�)�M�y�Ɂo�\8��&\��Cf�'����#�	f1=W��\��4�`�k�5�Pl�0�Y��D�`�j��Б�^IJ��!~HrT�d��D$�=��XZ�<�/�:x=����"�Ayc������۪��H�ޔƲ�:'OQ�gK�-&:��0u�I�Ǥ;�g��_�4"v�8@�� W�Ό���_r�]�g��ӎ�*Z	3�:���n�p�����_0��@���bq��:f��>��8��x�brڡ�� C�t/ �ʲ$j����WD��4?�V˦m����in���Ip��C�~��焤���D
���dg�pѦL \lW>�I��5a�;� �(��\�6F;ߣU��#�X�iػ��Ë�m�%�0��Kb��I�s�7G��G��@D�t�
��N��pb��M�=��b�O�`2;'�������(x����1J�R�Q�V�Q��q4�f����P�%�0��q��)�#�b40�v�9�8��x��ևC�9��e����Bf����Z�.��I���� Y⒩Jh���Ă	dT/�|@�U���	�1�Lπ��i�@�)o�y�YK���3r��Y���o����͖GL��1Wr}��A�����WQ��J%�l���S\U�kC~U�5��	�K���PD�u��ݥ3�6.2��u`��CVsgu�	�
b��x�;�"!u��e����H-����d��&�&8�,�5�G<%g�C?�����ᑮBS%�;���l��3��U�6h��z܇u!������톛��6qG?{�]i�7�GN�ul��k�z�%��
a��Q��B*�+��Y�f�*�Q�ȉh�Ӏ�1��X�z�UF6��_�����$t�"O�yYʄ��SBH�C5�Xw�,��='��0؉D�c	����Ĳ�֙�;���=l91h�AF4PJ9�v��C)���8!U�`G��������?󛨤'D��M�Nq�_foIP��5�0����h%�C�7	���C�D4�"�1Z����ɹ(h�.S��G]xZ�AH�eޗ�ʶ�[�d��!� ��p7��ߧ�"Mx��B�Q�f��ϛ�ؘ��i������_r�^�RV>�,`�fW̋8�n�����vѺ��L���V��Mi�/VWVo#�+=�0d�`N�����_.���?Pg�b:EΌ��[��LX��:�MU�8&�9��**�r�#"����c��_�u]6�S5"�?^2�4>ճ�7
#(\飧<G���\�B6��ځ���o��������?<�GiL~��"�C�  ���yTϵ\"���FK)˰����MɊ�̊m���2g����� /M��GX}ި~��|� M�;n��+qWC��}��*��r�����`ï���p���s	J�)6C1�1�"�����b�u�����Q�L䑄��y�Z�	��[�*,*��{gBU���>��d D���_Ӯ��3�1uVt�Κy-=e7X�^��xMƧe��|
�\��ᚙ�O���Ejy��b�Lkc&�t���-zC���'�nҌ�u���Ȫ��o+����3��y�4�Dh�W���rU��F'��T��Kg71� ���������Y�~�1��Cs��GF����u]F_�V�]�ǀw���4�Ԕ��sAW�\Z|m�K|Yԟ*_�O�#��u�6�j��QrO_=��Np/�$���7�oJ��e�W,���xϹ���,�J���0=�z2�eI�*]�+7K����ND6��̈Z٢-{��~T���~L���Ǔޓ�J��8QZ��8.�*��c�?ٶ�p/���m.�O4��N�����% �b�����4�+%�\��8�F����u�R�J�W��91S��̐�o���{��4�_D�䴝yq����J�@�[�щ�O���8�#ǵ�`������	;���f��,JM�3��.��ΐ�G"6����yǶ�<@� Ib�a]A��>v����6�l��TA";i��}��XI�
�T	�^��_�2��ڎ�t�I�z�_M����᥯o���[��g.�d���}����
5_�C�.�ب�{�K ��3F ����Dښ�4���6P�}
n�Zc��ٽjem���쓉���H�v����/8�=�;I�C~�Y�j�L���M}x�,4'�MVl����6!�H婻��0��X-.�c̶�/脂�ň�5���_tc.� �l�h!���5v�V�#�ڐ�Z������yW{��í�O�A.�̀��͊H����'�*S��D~ѝǖJ�<�NH��!Jt�Է6��G�t��AX
��@�3ֽ6�d�D"R] �3��cR'��k���b��|McyV�q�J�B\���dR`�[F����r���J|���@��;��K�Y� q�|����qA��2�a����*�+��&��g�NL������<"-�����n^���=�����Aj�Z�CА1�_�R����j�ќm����'��[���5�
!*�M�Q#�i�{�Xʹs�a84����I��H�p��I�9��Y��1�z��Ʊ[���֝�!�(��	��LG�=��J�+��w�@�U;,�pT�|8#à����J�Zy�UG�5+�"��|n�R�c��Y1'��Ǎ2��8:��������$ 4Zڨ�HU+.��������A�(����O�N_��z���QK���p��S���ˮ�H=X�$���C�o�7�y��U��ߡ0GM+GqV�AQ��������6:g�c�~
6�c&1SDh��Z�:T�3>8�]�^�rr6�kh�ڋ�#lK��%#t�[9#�Cp�Z^� ��[hk�}�eMt�I-�@���]6#�Z����@�)��	�S��#ȏcp-Y���{^=�$�矞�g�H�^�q�6H�ݥ������b ZD8�h}��h;׈_S�Z9t�},�Wd����QU�z�d��W���4x�m@��#_f�w&]=i�8+e'?W��j�Tw�@g���>�$�uA��ԼTpe�N�aF�h t(U7[ƹ[ 5�9����P/;���@�?��lTCL�Օ�*�1[��t���^����ʄm������_RLf
����92,�ے&�"vq]�K�����@Ѕ0u��_�W{�l�|B~5%e�V�� KHq�V�Q&�>�9w���Ŗ�:�g;6���1͊��ó|{�k�;�,%��#�܎B�;_���Ui�)��i�h�ߕqz��Ff��vn�%���pUH8�U��
[�kZ������&��x�
�P���v�x�~_�n)�v���p�M�O��	(�I�_Cw$��>�"jN`��Gk����vaZpCᰒӛ�|���Ξk�j,2xM�9�Vꤥ-�z�h��Vj)㱽,���!�lz����cC��� ʒFye��~���j�c��,o<ĺ�$����jqy:P5?ЋÊ�5d��틵�g��֦���%si�e��#g�yfF|�R��͌�d�І�� "��h�����n`^Fk9�Hخ�|J a����p�S�t��umv8��ȔP`���t��A�i�-%�\�; �/�����>���.��� Ť��_�A�&@�������'��"��c\9�5�l�9��3u�@�8�OW��W���9��/)SQ����>�%���æ���	��
<��]��c�@$�g��Z݃�~J�TS�MuS�P�>xhy��	L\G��>�m��Z��b�?Yb�EM؅���eԋ����V�4O���Дh�+}��,.r�=�9R�_A��Z�fA�.���;M_,=ڶ�^k����`>�L`�PeVw$B�V(8������4�yL�q�!d7=�XI�C�*5������c<Ot�ա���%�'	<��A�N��)�����y��Yv'�� [Y-�iD�(���#Vh���g�.e�),ؗ7hw@��H��5���B5[��o�䈗�v�+zј2rLٽ�Piު�R��r}	γ-&OU ���m;�w�noj�F�'5��oo�3�{�R��r!:Q�7M6�^��a;�D������t8$���`/=� 1�i�ʖ��t1r�c;���Шe�e�2/R �p{7�\�mD:e���=8�(�w���J��5�]8٣�-R	�OJad*6˰�IdO�:�g�,o���y��=?Q�~r��]_��mՖ,���%̃�������2��\�<{�=ď4�d_+��cݿ�y��<��&Z���VA]N	�J��GӅ�7H�������*t�Www�D
f�j���w|��b����_��3xtyp@w.\���I���Ni����jۈ��/����c�`O9h�>3�f���
���n�����#�j�)������"�d��6�NJ9m���M�W��Hh�������B�J��Z>ʢ�%���SI�u���c��=G�KdDђ+�S(���@bɊ�hf�TO��\��2:���b=һ��+��(��qx_�����F��|^���/��fkÃ��'?�����R�Oj�a{.D@�,b�V�E�[�1���po�qR�J�wF�Jn�h�kn� ��*K#H��q�$H��S7���o*�I0�v�d�ڤQУ�+�p��p����xA] 
R����֯������z����m���u�[V�[�1՚ƥv�Ea*&'�9@���=�F�o�/�=B@7�����Wo��7��6dk� �J�g��?�����2�Z?���x�t_���H��.����7��Q8�j����	���n�|5j,|�:�����_����'�D��mG�|������?oڝ���~�%���-�ޥ�Q�U�F>�V6�����@�ÚC�l-�����8%ZT���oLc�z��<jl��ڬ��ਏ�t�:�E�F���O&@�>���K���
�Y�����K��D�׸�
�qS���0P�܆���RD��ӭ����1����'�;#���-�����f'M/4���!��d�,���� �U����q[��(���D���,���޸��8��{��c���b�?ϻ<�ʜTZZ��I�j"Q,4����;���p~�+Q�wS@�3��r�Lx�@��y&)%:"��=�"���y�O;�2�~P(�J�mX��Ʈ�J0:I��3�]�^1�8��F1�"�h�u���!R����s�Fe�u�B^�i���j�PB���e]a�g� ���n;��wq���
��
���H�����r�В��
t�k��er����Dw܊��%��0�ǣ��͍(ne>�3`<����6m
@��4b��ᴎq֒ɋ���wN��A�����D�JN��=9�d��:PˏE�U=۶#�v�yii�_�{��dNV�-!����t5�v�T�_~~)y��%U�S�$p�(N`QA�Ua��s�(�A���!(�tGl�AgH�P�̊�$����Hz��jV|�Q*2�%
*i����A0�(;��꘷DHN�DP��vr���-�Т��	M�)��o_�$�Ig*dwrs��4��ao���A$�K�A��rLȅ�Ӻ�4<�m�z)�`~1g�>7R���SH�y;>Y�/fzu׭"������!Q�Y���iKV&�N�:2Ϟ+��J��j�[���)́D�o�3A�z��60��T)�*�bK��7�]�<X������i� �9k�O,�ـ�q��Īx}�����1����úhW,�^���������%ƕ����?� �s�ߢy8�a��b�m���,��֥̎!�[�?	��,g�t�����w*Q����lQK-+�����zL�f���g�9�p��844,vM�;m+��	���f��'Q�<�aH�����\	,2y��X��:$NI��[W��N�A��x���9�E��'Q7�s�ϡF��͢d�F�F��H�?|��ǂ�DR�gs���)�_�������������u�n-���)+��~�W�@q��ĝ�Z3%�S�>�����h�����z��Ss�[ui�w��h�Ql�$��П�g���t0�U%�WG�.j,��z�7[Ex�\�=`���.:�;C��s<T��ꦍ}��˼n����]��@�-�<�_be�̟�efb1��g���Xm$&��|�=�c�IAn�L1������j�xΉ�e�����"4�^��ز��;�ur�ZW/-�	��F�#���,����D�a_��$vm.x7�i��<F2d' �8�.�P��:�TָN:d�7��N�&��X��Ś���z�?&I9�qߎl���n	�;��L�NQ�%J���E�FL����I�E�i�<,;�O���/XjS��wj&q*y5����N���G��W`o���c�6.Y��&��o��ƌp���<"`�VfU-j�V/���,�1xX��1�]�0[����$������#�1N=�1f��9BCK���ŴJGG}���(*��=��*8��3�W�}��5˝��@�,዇c��5�6�+�n^��J�­-A6��d���|�䷟>�����e	�j*�Ad4JCe�����>c5闍�ׯ~�
!#��yb��StO'Ҟ�m8��L#s���y��<D��#�D0l�(EVx����.x: ��,���R��p�u��Q�	�Ƥ<I�/���4�?X���8���sߤ6�/����1�¢���~a�4�9����,QS�=h�G3�� �`�A��rB��q,�����aC_n2"ߙe5�J�bF��!V���Gv�'h�"���J�#��u�@�y|�5��m��Φ9%�C)Fۭe��e5�'Uw�`t�H�o(j�S1��yN�q�h%���ʢ�[G��O�c�0�����+zx�����>��I���w���`-}B��`��_��U�Xؓ�E��t��Ex��Κʂ�J�<鐠�����i��e�D�`�G���R�u3i�wOꕶ���gdɋ�z�łc%f��C��H��0�kͫ3U �����x�`�[�lFD��[I�6�}����п����ۦ���[pD��D03�{���`���-s0����#<;}�)�!�6����H�`��e��~������Y ���A\����Y��9p-����@J�(�oS�MD8�.1������F"��N�h�0_��D�^�r	��\��hLZ��W��4���������N����	��Br���,ӷ	���%��!�+@�Gr�ʵ�AH���[�C{���|X�y�X�C'�^�r�Ⱦ��F'|���K樏�W�x�k �n�=�/����-��3���/�x�T�y7y��e�y����na4T�����}@W*�]̫8��b7�j����yk���4�I'�j��26p��ƾǒ����*ޫp���hh�$V���#o�+�y�MR[mr�a!�5�n��t�ί:c�Aɀ�R��l��rR��ⴀ�1x���5f��RslZ��8�����mӟ��W&�� �����d�*�U5����&�m�|��B{�B�N������y>�n�/�Q׈#G����*r (J7��LVD�>�CJ�jL�I�X\ :KA�P��Jh�yP�sΉ" ��������)`kg��C���D��m�������%�)1rD����n1��A�[PG�3_X�	$J��|�av&g�k�Qt�d�C���eN�[��v���v�v2#'4R��e� x���p�W��"C�kX��VC=��o>[Սh����R�M(�R+�R��#�a\�i�;F�k��^ٜLi�r1Cե���2��p��Ռbx�9A�h�������:~Eې
n����eu@9���rX:kI]Y:tO�AU�:n�M���Z��u��I���Qꀶ_�u����3���!�"2Q���ZU��D0�rG��:}
�SDA:;a��7s����	�>]��X~"r�Tq.#��k:����/�{�����X�x�X�
� ���y-uH�V����,��*2cG�M� �&kZ�E�f�������᪔�KTLR��ղIz��L�*�,��*�h �&�dxWi��`Ӷ�keN����O���r�r�3���]/Pa�.;I�A��(
p�#*
��i�8�ϰR�( ��`iw��&�R�7�[���lRн-�67W#Ұ�	��e�'ӷa��Qu��-�h�y�V��j_�uSf�8d���ug\�o<��c�M�s�_�.����&MH#�%��u~�C���1z��	��%vg�6&5VQ�wvK�����FVr�upR"<�PMI������V����y�	~��Q������"���>��mJ�Eٶ�|8��2�=O�H�,\����J'�)�ӆD�{�kI��Y�C��O��F�T���j���M��`76�1�ʛ���3qA��[�g������R�7�G��ӵ�1FO�g{��$��·�eT�a�i?���uZ?4���ѿ�A��dhмm����ۆ�"�7����	�amx��������M��Ð���ٰd[i��wL7��E����Nn�����cw����f�Cl3
�dPy_Vӓ�z�&�:I�N�D�h����Fs��|��q�u�|�n�6 ���%N��0&�� ���@;׆{�^n�rH#�a)]_]��	�FX[���V��ߐL����͔����$����K�b����ߗ��A�����wShYX08���_�`���RP�b{����a7�؊�=��k��CÀ+/s��(ȗZ	���\���S¬-�Z�����OG凝���Lx����ven�/#�8�Vف.Ͳ���s���̧����}�POfŅ�$�	��>&����AUksE6֨K{	'_���$�0�+�ҩ�{�yj�K�ZH& U��,��VK�7��1a��jY�U�X�J�B���D��p%e_�7یJ����.mh6���<��s�"N��A�;��c�E�v��Y"�p5	���"���o�Ĕ���#>79zĄw�˵6���;&���	�����2���L���$��C�)#����]̔�m+����2C�ϬGޙ_�e���,m�ٍ�6�6�� c��kO6�ƽ��*Ɠ�?R�?� +z�Z�I���L��[0�l�/��c��4�#Kl�J�I�q����5��sF@`�nT-�=
�m�Cc $���P�6w�v�����Q�ކg_��Z.|�nh��'Fv�H[)L�Vd��i5�ŕ���v�8�@��"���ZT<%�ڶW�l��cz��M�w���g�ع�_����6�'��Z�����a��.���C�T�i�	+w�V"L)�����0��Mh�S�q�Š�_��gl|I��1�($���m+wJ�$��u�w.JdM�.��&z/�Mh0%�ah�p���/�e�ܤ���/H�N[$d^G)�	��z�+q'Xm:Y�~tJ��nE���lzX�l%�/_E@R0?�C�u���>�a���i������
i�0�*?S�6���Z�l9uRJ����0H)9b��� �"���t���]��S�nN�p�'�0LEr��V����)(�Z��F?�p��!/M�`�nD�鼷�Ԁ#4��8{��)
�I��X��e
;�1QT�Ah�zo��M	���_��\㯤��3�rq_bӛ�����Z�L��UWi�n��ȵ����p��{s��D�}8��^�5��Ɗ�7V��D`ҵB^���;u}0?7[��we���[s<�T��0;9�l�+����Nf���&z�G�}�V�N֌�o�6����2�J�wtVD�o,�p ���}1�ݱjNP���J�	M��S\�pˋ��<i/s�����f\s��K���χ�ʡ���I&�>cB��:K �s��Ey��x�/��)b���J���~����kΞ��շ��(ie	�o��gI>G?U9��V�be^|�cE$.	
�!���F3���d�d�: 6E�A���O�`�d�r��K��y	B���IU+�:~��ĩ=� W��LUM}9��Ԕʢ���\�h|�^WP�1���Y�*[�ы��I�����s�BH���#���
2+�zåH�Д�4=���gb�.�;a챍p���m8�6��_񶯰��";�E!T�p�pi�z���r����
G�z��֕�B�1|\B|:���3�9٨M�f��j����m��G� �q�wJH蔄3�f�L�ʌ���o�m�c�f�q�wY�7ފzQc�'�>��3�(͢n[�WE����`�ɗ�d�B���B�˴u�	e_��y�4![����}2�_�Q�k/QV���\��2 +�LZכ�yL�К�5�M:�Qf,�;�q�,X�QuB�v>Ӹ�;��d&. O�w$U��X��-�p�GK1�C�L�-Y�h�����Άr:�ŧ�S�'l�ŰTO�];-s�b��z�Xj��н���'�3�Z�أ�4���k�=�.<a#�bYn�f��u��'��x��'Z��DG�9@!s�(�_� 6�p�=�{�i��~���]{�IJ.{����^i����V �~xf��ތ@�t��x�X����L�S�'loZV�),`$q`��W��P"�(��hGO���y��|2�ȄS��J��ki�>,�8���YVz^���EN�S��	;��ޛ>��OΗHz�	Ɂ&Ab޽�D�)8/f�)h��]��\m����A���	�)\w���du�Pߑ��P��D71��F�hg�}�W��$�����I��#@��˼Ґ��h�8��A�VϹ���i4���6��=HC��=�ۣP"Z�cJ��b]��=S�5��,�n�0�4�g�DX�ۍE�� 1�!�Y&��
�2ay��KTl�'_�����[��N��5.�R��1l�D�8+;-�l���o���Ͽ"���lQ��gۂ��t<.	8x���I��`:B'�mM���f��A3��~���8�L/Z���4�O� g���0�,�?��L������R"oE�)��;;��g�c*��qͣ��|DB~}0��>���x֒�o룧�.7��vNa��r�z*8ڬ[��?�_a~_�펰5��W/� �H��0L-^���y]#�|cW�[s�_��܈����ӹ�^մ�D-:�׵��I��	�n�Xb�%)�$d��>��(޿a����k@��*�1D��2��A�>�k��$���4<���f��$�X��4ȩ�d��TS��㑩�qJ���8)�7���M�O\g�&ʉY�)ΫM#�V� `�h�#VNS�-HP�:����&��t����\�2|��Z*�����,$��7��]}���(_8Z>6b>��S�p'��3�5�!L{52�?������ �kg�wyk���F}���H*~��H�@X���?�L�7a9�k1v��\�);,�ɮ�1*�c�R�}�m��Nd8����r~�E�H@龔�('�6��~���� !V$�����cs�@7�Qeh�j��(��S�1WP�S\�~NK;��� N�>��z��wx����V�9��m��a�4S%�,m�@�9�AU�Τ%Üjrz]��P]s��ۇw�����d�ݲ$Y���/�[�t���:�%�wo����[���� o$��`�ݻ'�4!�?�Y��U��;n廙M�ô����i�ꆊ���� /�)9��t�H#(��6'���G���~�)[����iFT�3�sw�f���-Iym����p��[�N9EkƉ���������C���5i$���/#W�Kl��j�$T l�O)�PQi��S:~���j�S@�B�%�A�3�"��S��z�����p0}l{��7ǐΪ�p��Yl��e��>R���Ik�O�1�0�|={���X �y1��rv'�ఇӆ��XQ��C$D���6d<g!�d�0(���Gq�2���۹I��D$�(���T|CvcL��pYF"�2���f�f�������/��_$ŋ���t$׍oR�Vrq��~`�m-^�e�@�X�a&Q��@xPwS��7�ڟJ{�l�X�aZ#p����W�п����'�i��
�)r8���#�("#y����A	�q�K��H��Ü�sRч(;��R�2�w���b�m��&�%��h
��qu	�HC~���`*��߯[�	~��7���ǁJ����;�f)��Z��d�����ɉ���ދ6�Çܕɨ(��.��o����W��=r(��k�B��D����`e�u,}~����TJd�v��f��;�74��ZXj���
��
�H搩�ۍ�k�;�.��A7����V��?�@��>�2>�Eg|4�Q��qɛ��=Ȩ�&0D���h������Q`�fԀU��,��=i�Q�a*&ɩ�w���sP�9��+��χ�e�K����)��m�ZM���t��h��spX>�r�B��D������f[����3}=!1�&�Y* a%�SN_m���6�kҐH�s��qB9wb����y���g � ��>�[����9q�v�2��N�Ǹv�	�K��w0���W9�c_#Jl
e�,G?�`�]G"�CJ2�L�,��rb��~n��(��~}��;���k%��B؇����ޕV߈�ܤ�qڏ@�K/��)���DE��D�;R��Id~N��M+�,���،a-S�
�L�N��)��x��ɼ�FR,��;����9	@�>�S1�H��&�t62�a�	�7&7�t���^Q�����6��+>y<=�:zٯ���G̶��q?{N0�;�@����T	�~���Dī{���W����U��� �p��h��e�uޕ��;�:Ab�þ�u�����`����6{s[�^g{?��8�l�X�D�W����������
C��E��c"�(~|�K�� �({��~�M0��
�[�
X�MH?PW'oZ�q �"�2������9nrlx;�<��:R)�@VW�2>V����ۚ��
ޘ�dR����7?je8���Q�A�Î���g� b�2dV��Z��@��_�9~����XǗA��q�&cA۲���"T	?\��ˮ������<��6��R�λ�E��v6�l}ꛉ��!M?`S��*A�]OC�K�$�O��:�V<T�FS��_<w�-�84�h��x�Ȉ�����xP�h�>OW�m �l��\,��O�qS���7�o�t�6�!�l����VK'4?�d�����[���S�_'��7zw��ݟD����ӄ;ʭ0^�]�qk�~�a���r��S��~ܞyY���;H��o�ev:���6�㬃[1��?{Ӣ�r��Ĺ�vj�N񚣜��0l@#|��l��0}����Њ?���,k�vFuԴC�
�^�4j�2��.����M������4���V���̜������6Q�n��K1-�Q��4T�E�~7&�S���x�$�X�Q��Fy$��B~��N���/5�u�K2!��G�e�g-����o��W"�a�>�����!�����J�sz+�\Ѝ�_�
h]�M$خ�?1�|R��]�"L;��9l���6����-HyK�D4�g��*������!ж��/*$��0�SpQ�]0�ՖL�!�>�{�����NW�j�mA�%�&��ڜ�}WĭWf�Wn��r���2�>��E_O�����LZ���Ct�(nn������$��5��w��C�
!/T���_��H���5%�$v�/w6v)v<Otan��m$��m`��P����ZR�@cP��Q���+�4����^ԑ�]��IF�^���@|�K�J��3��P�R�r�c����5^L���'O�e�/��цK�k&ç{�F�����P[ڼ-�)v<K���ůz��Ll�~���*�"b���L�GHŉ��i����v5m�ϧo��8_�v�(�w:�S��:m��H_����Tĩ�{����"4ġG?<�V@;��.+�Y��	x;M!}G)�;��e��ۯ.��Q[!:�d] ���6z����0�N�w�E�ѱ���;�Ң�1I��30�v�{歱���!���#�r�w��h���R)��jЉ�/�5M�bNR���u|��W0�����=:KW�Dp�����A���|�o�������>��D���]��U	�P�,�Ӟk#���=�A��)aDȬ�8!��oơ4�ggpu�a�^T���S��xb�vY!��>E��Z1��~H�>e���RA�GC�x��UMX����4$Z�U�����H ��/s��{�����������}?�!���-x*���mf��Ґ�F�a`�#b�Pw�}�9ʩX��w�k��Ҙ����3�g5��+/��B���h��m�7o�f!hr�<�G���A3̶�;�`N	��u^�D{��w}|߈)�4o�� X�HY��� Ϗ�o	[N��ѩ��PIe�5��?a�S_r���9�C�T#���B�U<�gNO>���%�e��q��º<ɔɢ�2ز2�djS/�-ߎ9X!� ��&$�2gnL�9hT�1#�/v�`��L��p_ ��'LY�PU�]��/)��BE���V&zhOsML�w����!I���G�W2���-ܱ<�|����}��k��t�;��U�Dؗs��رr��('0��D�Q���ۂ���5K{cd.�ܵ���ك��H�Z�{{y��n ���G$|��`��z��GB{���0y�'b�LK�v���{k�f�1���a�ņ��i�|���v�U�M?hgg���)�	�B�5�o�r	z7*����"������i���_�W�9�!T�4���d��$�P*M#��o/ϋkInD4z�M,�餀O�1�$�J��+��~���I��1�o��[Y��\�b12ɈUo�E����U��0�8̼m�44?$d,�� <�I[��"t��q�s'�-jy'��e�L�RO�>�����-UU\fֿ������6=/h0�s)��s�c��z�D[�Dح�e��D�* l�V#dN��|{��;�kO��r ����o�[M�B��""�5��~���Od��
�}���˓������A���JW��O"e�1r���c.v#�l_12<�#(��:L��d-Y�6�o��P:.(�0��n�9���D�N���:�Q��P���rC٣�[4��cΆإ�5��s^���a[㰕z8��*Ǜ��+��~ӵ�x�Ceu���-������خ�Z0��q�9���=<����^�u�j�ٙ+�ߜ��s���+�h��v�}���Xj hu�ȳ������I�AՅ]�8\��c��/^$La���'$U��qi�c��������(��5,�9�~0F��A�ƹ�,d�-�ԭ])q<��#(�	^�ق�
�ȉ��F���0��`-a.%�~Y�hc�0/�h�G[")��Ϩ���d�8��Ƨ:�d�A��a�=�b�9ܻh���{����""L0��l���K̴���|����^�W�f�i�6ϥ@L���,V�Q5j��I�@�J�����бD�M�Dt�g�����~�P(!a�r4Y_H�y2��A$�v\�?�ׁؓ��+��XhiU/ ��y\ödA-������
�z2�7�`c wΕ⃳
↪�������p%�D�T2(L[��bΰF+y�95=� 
g��QG��8���sƕ������j�҈i��N�#?�}��J�d-�9EH��ė��,�������b�a�^J���Q������И����Fw7���3��	��{�/�w\���G`������<==��Ra0�ط~ϥ}�)�{�̈�YW�D��K(q��v/�6�uT���;*�2}���ν�$�Y3pv瀌�H��V�l�{s7�������2iΚ�������Kf��Y��Ju��ժ
5�����e��Uo���h��ȉ�k��)#)�q����P	�>�D"p�T� �9#$�V��1��7��\3��_�Bs�U{�c:ꘞC(�$x�� ��uY�4m�PK�nF�K�+�������5Q9��f �����'��_��G�b兕--��e��Ȁz�����#��ȣ�Ƴ��p���<0l�o^ܖ��:�%sG��2�D��-},�+�䐶ESe����H��[9Fr�Gm-��Bl4���5�Ѩ��_?и���m�I?ۆ�}�
ơ��S%��DV��֝V�	ꏼH3f��l^T�QkJ��0��3�,[�+��[�Mr�<9�~����:Hg	�13NFI	i�ը�u�bp��@I��V��k�/tm35\�����\o�2j3|0�ﱎ-=ap���QщXb���}G��XG��*5������	Go�}��ߏ��<�{F���Cσ[��E��23?���q��SpU&L;�5�}��������6]NHw6�1�PY:�{)��Zc��Y��A�e喘�g�UP�]��fG�D��5�z�"���q��H�6t�HM��)�tv�ғ�"�K}&��C!Ӊ&?�I�?�)	�M�QYcS��'�s����Z�|�C@��5�l)n4Չ�q�dl[��A�����;�;���l6!���s�K��8A�T���)��d�B�׶������M/Z�5�ؠp�^y
v�;�!�����;h���[���͐;�=�i�M�;�B���}�I�b�Θe�7��VV�Ci1��Ժ�,p���DǟH'����/#�T�Ρ#ȸ��5U4�Y`E�.hO�d�K
 !)əd�Ƌ{rI�>�$���)��p\G�yVrV����)`Q�+�*����\5�8�yCy|0��$���N���ݧ���_��Y�5s��j1�8���6*�K�����F��h���KSW�Y����v�ݎm>hH?���u��/#X{X;&��R<4�f�S���hLF	x�)�&�Ɉ�ȉ+ô��K�������o3S(E3�E'< [��=�{���T�%]h��MF^E����d�u.�4Tp81�9�hyD�K��3Ղ�6Nq�d폫X�\)��f.g~=z#��}G�'����B�\tl�d<����>2F6���r_��d񽕆���ڥQsVxb����nت��3���Z�>	T�8���E'��Q�>�u��x�99���ѯP�<	��t�{WJ3���;K0���Ʀ�&��3������zG��ѝ}=z*�F�+�.k����[�e�Ҙ��%�t��|����Ȋ�k�I讀�V�ϫ5���[������֑1��w!�s��4O�������Θ�YѤ96h�aM�H�g(M{�I%~���� �[Y�F�wY0SRs�M~uvee�s�V`ʈ�j���_���:��Y��(r�И_	��ϥ����5��dupy#��G(u3 σ��2�*��\���w�B�����<qJ��l_1"e_�xiA�� <uyW=y�2c3�W\�i���XO��A���\�4d݇[{_����9e��7��46�Y� /�n�#�>9��~M �ا���?�{LZˢ�Z[�H٩
� 41~��D)����5�	�b,
Z��寀�f𖮆�\/��
`I.w��cy5C�E�!4���6/B��߮���5?�� Ͳ���p�\�:TV/�[��V#�͌H'�;�d��:���F�Ѿ��es�"��	�D�j��Ӟj�[�i���xt�3|�.��G9���wtU@Z����xC�M����U׵^�K��7���R)X��;x1�T��%�UR�gxs�fa�΀�rBs�a��N��W�����:�J�uĦ���I䜓_�,[�5ov{�t�����IMCk��RC��d��7�h�|���R�0�4�2<�K3��ųm�B�D��Q��)G����3L���hO,��ע�K卥��a�����k\*e[��̃��7��ĵV�;�h?oa3~�f|���$k����U�b`dA�VZ�	� ��)~�`ݐ���|Z�����K���MP^�Z'TD_RN:�^U)'��L�S/6�8�~�P��n�/GI`�g���__�F̣�ڬ)*��S�i�SKW��=��Mj��/�o��(F������� �S現�?�s��n���(���(Oo.%�4�e��a��_��������ʐv���N{��M�I`�G�w��`)1���0K�`Tf_ͼ�W��wz�����#~TOfi�R���������Vr��´��g�$
>�[?��p6wa��]�ˏWWZàJ� GX�"��������-�c�ͼ6�Ƈ��m`����ΰ������S0�;�u5_�d���!�X��})�
4e>5R���CN���&~��ɯz�)ْs̷[׍>�T�pyL���Da��F�g>�}�fl$�FG0�W��<HTW.�[��T� ���3���!���f	�dR~H�8�)	��i\�=B� �^Gq�N}=�"�vaH�w�*�f?���$�aV�U��imC�~�2�h�
��Y�&�XJ�D��S����B� �J�q�4��<�3OQ����^�2��J�3��3����ȁ~�ڱ����&/�B��%��9�u��'��ΐ3�\Hw���-������6a^K��.t;uv��j5;�Ҷ=��cH�S��C�%�w=�;��X����>�0��:fF���KaW��8���'� �\M�챵�i��y��]�����N||1$YЈ�'�R���P/���Q�[���/a��o\ԑI��&���Ҿ�6�c���������'A@l(���g�ɮ(p����g�@�D�:�4�.�>c�dU+#����ⳙF*/�����xԧB�#���W2h���p\ph��0�$� �����O+b��W�[��&(���=�����e��^>M������S��7/���n��Ur���y#��#JvX�����̾��Z��o�E�9�L�]�A��H�����	e�u�VEr
Z�f�*�&Ǜ�8��E	�p���� ,�iA\ea�r0�`z��s	<���#`�/�.�H�M(�֚=ѾcJr3h�(3�Ƈ"�=�&$&I������8�;>!���+����G��j/�r���Nm��*��1��I/�dLSF��U��]�VQ~�r"8�fˈ�������(l��(D]`?B�7���\��C#�lW��YG���y���,\�r`Ww˅.R�k{�J�1d�/Y#!�zǅ�w�ߒ�N�#�����!�_��q^��k�dҺ�D�6�ǂ{�M��hb�U����) �y'�J�f���A�����L�P�֨�NV�g��k&��T�"�/��i���J�Iw�F�U؏�g��N�	&QGn\|�����nd� ��6�v�Oѡ�R{�W��aߏ��h��l�ò<z7��}�H�:\�|��hc�����J��e�Z7�?�HU.IG�Vy4P4[I���&f����Ȥ�w,C���猈�i�}�'D��a��Bɴ��d�N|:Î��Qf�V)�����2JK��O���]<XL��a�?F���um�p
�(/�S�I�,<���@ �0���f9'�uᰘ���)��&%X�rsk���?K��Sv7~��M¢��3��l�Wn��g��5�ÁS�3�o^��vzR��iǙ	�²T���\W�+��Z4ҳH�z�)�]5�ӎ����XO��i���|<v���=�����OEZ��_�_�C��������Ů����#�bt�l�6�p鵖?�E���pйl�;p��[�HSR���N������`�ֵpVTjC�=�`ʺK�D��{u$�O��b-�V.�qmzxb�i�KH>��H���}b /m}D!n:j��*^��?^k� ��k*�AÍv+Mv�E������|�H�����m�L%�l�;5F�tȉUzGL<������uM�	��A��'Ũ�º}V��NM��h��p��{嘊�E�*j��A9��ΈVGh8]WhЍ�`�WLM��\�q��n��W�7�ou�-�Ͼ�Q��.��d]Qn!=O�u���I��D�O�Cl��0���H/��8�˜�"�L�*�ۉ�B2�a�B�l�p9xDo��4a{JoJTJ(�̪���� ݧ�'P��]GX.Va���nB�R�ܔ��*�i�R��1TE��X���h���w̶�@��Ģ%Z �� ���1����-e=��`"F�1zؖ������ۓ�����/��G��1���&���$;ggb{|�˸ۨc�]�0f�=�.o����0��I�N�0�[�St"�K�Q�/�ש��87�w"jK$E�c�ě:� U�H��XU6U�j[�r.]P�ՉsO) ik �����/.�u����O74\h�9p��&9	 �/6
��d8��=;��Ϥ�G��%�$P~��t�;��IŰ.#"��n��_'�E-�����h�*9k\�	�Sv �K�%Ui|/�A�2
�H���ekL[�>_-k�?w;J`݉�.и�=���[mR�CN�p����$�Ҟ�BQ�X����2�&A�H�Ͽ6�}b�u������^�ѿ˴o��ڀ��ᶽ/$�� W�.�Fg�*9�o��!mj��3?�S�M�	W%��.����5�oU~{��@��
���^�Ku�7�v����`��CI��<1/k�WÛ���1�����9������I{͂�S���Y�c�uh��r9-�q��.�گ3���-
g2H���K��k#��.WA�cТ�Nu��{CRq:���M m��X�Jȕ����Һ!O�j���t80��&�EB��fӎ&���=G<���	�y��
�8/�_�4^���['��p[#��7���y�����)6������Ya�u�p���4�����ˣ��O�Gg����D%$u7Vcb�(_�!kW}z��䙱B3Z�BV�Z����׾��?[	8hc�%�\���7[M���3�V��.�gP��QS��`�Y�1%=`xO�����5�B{2����I�^2#�J/��֘L��`q� 6�x��+�������I�kS���C�S��^������\UL�=:�����o���1��׮[�n��l��p����������p~S���3x2����e��NÖ�,w���d��������V&!�����|�E�u�C���W��ǰv�1'�D4__;�lp�^y�7����U�r�7?��!����7X��g�q�A��Tף8�5I�:�3c� 3S�f#����͡���z�"���2F�XO��L~�z
��9`�H�I���o��8���M;ӒI�-��uࣛFYQ�Q8I�38>Vգh���\�<"r��oJ4��i��<���E�u˭́Q8y�A4-�yU3M�o����B4�C�K|���k9-�YYn뇌=�LſAz����ء:�WK�R+UO�F4��n2O'`r7p���',&����P�0��ȫT�i�B���F��Z=���ؒ�)��d�C�ǆ�����m~b��l�w,U��0Ͽ$HH�OD"���6�6����9A��y���1��b􅍓��5�R���;K�=�?p� �4�l�y�rP���;��'�ø��Z�o��b����"0j�-�s��}$�׍��dd�8B���ⲃ�eS�_ݰtf�Vm�\��
��`�@˯?���5��y"��k��Zu{x�Q[�n�/�YA2D�ff�V�&�1]#��R"�z���ܒV@s�nsԻl�����Yk����gp�������~I|�z�mDu"<l5��_��W[E�<~i�^����T����o������4 ͿC��8�,8���"��Sj�b$�&iV��J�M�~3K��S�
��Q!�ێ<Ih(M�uB�w��X䑎�n1��A����+~۾���k�<�G'�獷��&�2T�i�����ѣ�q'�W��j&VQe�.��Z�w�g�Ƴ�V0�2OHd�4^4�\��A�ɦ��§�%_��d��� �Y;͌��>2�œd��a�bv�
�8�!������-���鎮��W�h�I{|?�/����՚!:��u����+�ݫ���h���MZJ�d
�Bc��p��E����IN��~)0�m��۟9�2��W�,�}0�$V��a�jg���T�f1���1R�?�|�Q��[w��ܭ�����j���I�oF��f�ۍeM�i#ʶm����⥢�G��|lz���B���14���[�^���0�[�J`�*ϚK��ʎ�����D�=� �wU]m�eJH�t���݀)r�Bɵ�0��I�{w�*��E�lt\�t>��̽��;<�a�Fg��a�SE��h˺:��ù�B�M�3���:��U��F_#0ʰ�`M>���E��'�=��.o�ϸ�>v��V#�N.Ų[����͆��r?��F��g�sJo�}�o����M�~�;��E�I0\�1Bc���=7�ޜ�׻݈����&o��dS�hu�v������[�D����4��	K 'I�?��_(�Q/�)�4r>�`�
>��0EB}qV0��a b�j��g��\�w���O�q���D�A�4��c�^����{݋_�-���ל�C�S��i��x��X#�(��/+�[�!ޕ��-i����ǏFG:	X�������l��	O��c5U������z�uț���>gv��*���f���t�,��s�L*#e]p�Q\瑋\��({����X�|�a���q��XZ�k�$+��SC5US�A�X�c���K��M2���D���ҢM!��̄�]Sj�cQ����;���"S?3�=���V$��8'��B�g����Xsiv�z�����<Ż��s�́5
���!�����C�蛻��>�h���l��r;�M�1��a�����U+P0t�ή�x����Z����a���yI72˲��ԏ�U`إ�{\�#lSݑX�Ϧ��l��|)����z�_0Q[:Ï��b��@L�eT�6��|��x�{��R��H ȡJ;�^:%��-�w�Ru��=��w�X�6|b��L���w���]Z��ߣ\�Ǜk�����`)��c���jy��}r�1���-i̳��Ԗ�7a� ��\W&w�h��͖��$�hÚr�JT���Msu�O&"�	��Y-��<���%���/2���H:)o�x�#��nR ��S���]+��Mux/��L�$W:��2O�\Go�>6�� X��$i#0�o�z�.�@��C��5Vbٻ���3�sFL��o�{UE���!���T5.ʤ{�I��f�J�bۆ��^���#�Nw��a[�.G%��s��?���g��N��W�l� ���X�������J���㨊�j29鸈�$���.�5�{��Q�D��~��.�y 5��o�s����Z�"�?����&��v�)�q�?P5���e�8��Q(�	�-�Ko�`��t���~�$hE�ҍ�� D�����i�^򼱜���w�P����������Z���H�B��a��(:-�~�KB+��Sq(���G:b�xL���ΕF��Z�-�-����ִ�N�)���ްM&6����߾�05VA�T�ʚR�=�ur0#�ײ���R�q!���"(�D,�jȖ>���њw�AL6[+��H�����n'�o���N���L	�%��ͬ6�º���m���<��af�0���>t���/^PS�Y�?W-)�i�"I��#�Rj�$�G��q��D�h�O���,,4�g=��:j=�-��87@bls�.{�#M�a��,�6��>��L̙�&�QrW[��N�9�$#�����9]��ZMd-��\�W �xCB�Yn�~c�.�/I��W�]���3�*�i@�s�	+�o1��U�M����q�J3L0����;Z� ����&@<,S��[��&�Q.("UDvds �^"�޲*��p9럦O+g��	̐ÃDxv=�<�l�I�7a>���T�̊T!�<r2�g�xj���ګ�;~�ƹF�
�U:��&�h`)1t��3Kv��Ġ5���56��!��TJc%��'=aKO�~�����>��ǵCDb�k!�Ύ��5Qj=ƛ�'g�W��O(,���A��Tn�$J��H/#�Y����Ud+�!fģ47�Y�K	.���y���Y?7�iޯ��.�B'U���U*�|�cv`�F'�r8�x���p���R\��}�I�k���B�����s�;nQ��J���J�)��A[�J'c_��������&�	釖�-ʁ.�0~wY�b"������P�o��O@t�M�<C�x)VqE^��u:����
"p(�~}�b*;3�Jݔz,vA8@UB��������Wm��419*y��x��s�C|��#x�ETS ��T�#h@+��f�BI(+$Xyk{t�g�u<�$�h�n��r)�R��M�:�@�~l�ĳ?�BZ?�����u=�f��19�?��R>�dC���g��ox���tm�7�?\����Cߑ@����R�����IvM����(�m�7n� B΄#'���5���P�yFA���M��S$���O=�>�{T<%�d�3b��
gkfpRAD���ti�w��,��<�9�u�B��2
���P~2����R	��7�8~e�ɧ�z�*�R�8�73ꘈIR����j/�$>c��ފ9~�L��!���R�{������Rq^�{$���=�e²-�e�i�����B��0n;�-L�*b?�b�<|F���k�!�&1W�kdv�ɺ����;)�����\�=�P�遅����ݕ�`h:�2��?֥%Z:s�#ʊ��I!·��)f;�z�e=i��J	M��N0��@c�Ԅ9s$���f{�-���qe[?O�z�֣���ޯF��여���x�F�/$Y��3-0����v��*���#Rӹ��]��S��hF�� }
E��<:㈣�>��0���{16/Rّ�EV{��S�#���Ǚ.� �_��a'";���'���`�v�ϴ�`FN0z)h �J"6wzZj{�< ����mxT+� U -}�$d;����U�k���vuk�࢘[?��&���Q8���K:���%Z�k9f�t�H���当�ͯD��Q&�z�7��B��1�:�&��;ˁ���Pt�c�Oۢ6��&��0P�����9-ٵ�e����K%�i����(��Pg#Z�Z�;�����Yq*kt��p�'Ne�z,re��9���wӪ�Ρ=��f�ۗ�z��8��Jwj(����ZΛ�_�F��e��~���2~�t�@*�>�I�|�(<̺%���l�s`'� Ǧ��k�����WD�̴16��@�,S=?E�z��iu������6� m���)��!+B�O��y7��tR�����"����ҩD�������?�r[oƔ���Fۖ�����b�e!�<�5��W5}cC3�Y�R�i���qf�'q7�M�a��]8�:��9,>��W��a)g|��!՜!BO�:��N��1�@Y�����ű\�Q�����r"���Uґ['�a��Z���uF�囿�S�A�D��2Po�����GQ�ю�a�?r��/m٣�b3�r��փ��sUO��7v���L������V�(0���p����t����H����h�t�W�15��$�K�s��d����Ah�]x������HZo��X�I昖�/�Y!�\�'u:�����+��s�$V���ϛ��
O���c�N~�-�2[�������-z%���?���خ�/t�]���qaX��&��푶2��t�Yx�1���R�:��:N��L'��צ-o�@��>,PmK�� .5���a����;
��-&s[�$�uV^G@�Z��B_`�q.���p�i\/�*=�SI���>
����z�kSv��eHo�잸�^S���ͱ��6����Z����a�
�YQ��=�� ���!��K��T�%ސJ�b����pA����v��*?`]a*�>��"��O�����P�4�t�T2!��1��%=��J.:^=a��0���<��|�Rɽ�>x���ڡ8�Ȥ���������;%yO��TZ0�TT���}� ���WQw�9 ���q���16�\��|�P�[�l,�|`�k� ���<MS1���7�5f�]Z���4^�p$���E���i�^�^Z��6&���T��e�O�>���H^~������ �0�؃O�/ܵ�IA��/!޻
��k�3]�7����:e����j��ZjR��;��e}�A_F�Z��ל4�t��������H�\��x�l%�̝��Tj�����u��=�3�̥�{l����|�ךF
2�)$�����c�yE7�A��|�.G,M�U�E*��k�hQ�Vw�]���2cdka�@>� Y{��j�ys�I��m�;c��>6����B$t�@��6���Q�Asa��Q:�1j�Y��(G�s���²�ζ�v���w����g�xw�bE?A ��(d�}YgY�!E��P\u%*�����E��9���J15_�l|,�����ˁ_�8,F �JfJ��Ef�����Њ�����/�&�8 �ʣ�A�:�@,<�}����i�[v]��;�Q��0��}`��jO���d���7��'xNH�@z���-�����㻨�3��@d}����G<��f��X�) ��t�!�e���1��$AX)H0��� �'����{�aD�������I���cc�dy��n6?u�O����(�|���,!���9ʴvˢ�M©����� �^TX���  9Ah�ϥ��c���Z�);�zF�{�n<I�s3�D��2�ӧoE��]�[��֠`Pͳ`�8X`���ݳ�?!	G5�n��G}N�|�H��۹�XX?,�؜s�h��.��p9Y\�e:� ]EC�LR@���>�Ͽ��7��1��,��7xʖ�a�G���kA�23���W���e�;X�AjK%�bN�-�ꌝZ���E�*F��8v�� a�����l���U� T*.���v�gǩp}�P�O�@�x��EC	[*�'��`9Z��},t��x1f�BD�0	���D�~�`L�����EX|��ٓg��5���Z�z�θ�X���E��Ĺ����ՠ�qx�
gX8�3��{�K�H*�	�y(E[�{����x��@���D��O��ը=`y9ߤ�^|�f���l�z!���,K�Ja�"u�yim\`*VlGjQ����ν�W(� ��v�ͮZ��L桛*bP��mB V�3m	�b��:ï7�C:�"�$0���p؆
T4,�^g�~D���G�~���cv��4k����,�l��M��)�Ly�Ӡ��Sj
%b�',�1�x!��f$d6T`l��-�����=�,�ϖ��M^�ΐ�� �Œv�5��_�Q
]',�p�	�	ݡ��^6�3V���w�w��������*2�켨���A����]u;���x,C��X�~<��*�H[�=��+�r&� A�q�t��x�j8I�Q��u\�vE�K]g�	\���0���e2o�X��;�d*�w��=�����첰Ǚ��?	;J\�������I��*��%̜�@`��\sA?��qJ`!�x�D�0��y��u�s�:[�mK������)��1:������ ��n���葤�=���k �}ր׃B� X�V���Tr7dC�&�N,I�&�˳|JE�]j���h��e�.���j��.���Q�_������iA���F�����J���2�9׬�}r���ǀ:�l�3J��-@	��;׊��k��r�� ��N�&���.�Ҁ4�]�&�jW���.e����[O!{V��_yK�����iY�#�!�V�@bU#�U�^����P����w�jg&��h6A ��0\�U.j�����A����]N,
�tm^��s�h���s����n��1+>��DA�}n��G�)(jǪ��Q &�Vv�i�te5�H��F��ٮ�<$�3j�y9QD�B+�H���]�ل
�Քt+��ۄh�N���{R�X84%������0���l��	�ePJ�D v�i��Z!����Q��H����h(��7���<��އ�9>K0�I��x@e�h� S�rFz)u<K̕�c�Hb�F�V���k��C]�_��^�s���c_&�H����ւ}/E�x(C��dV8[(o9�����!��U#瞦5[�͓c2z$1���s�՗��B�G�Ƨ���y�Y���l#@k��e����������1�r�꿖a7!�� �c+�T��&1|v�OW��`�Gj���a��oa�� ���5P<�>�x��� mUϫ�?���s���q~�S��̳?Zs�	�=��.���T�b���M6�۫)��Y�u�4�M=�L3F
�oQ�I{�un|��:�#�3��"rr��?5>�%pQ�%_$8���4�*�W�Q��^I�+B_�g81��y��,Ў�mMTSg�5��q���{��&��5@�i�DSU�l���d+�l�_v$A(Bm!o��FF0HWb�e~���13Ӟl�?�R�K�P��8u�b|F+)ተ6���LҦf�^�9��0�3�����<K��������}(ɚc��p�/�f#+G��W�\� �i�-xjHg2�Uy�o���U���]�-�.����c��`��9��ޢo#]>��}�9���E�ɬh�V��]��I5L�!�U�O��hkF��%0��ݶ��l˂@�	�<o�8�t�j�(��[}e(h���K��3�vP�wg��J�X�Ɉc�_����H�H-}�~QR��c�G��;����-4�͈!�N�^��V��o�� t5�^4%�rnO��弓=_7$�~�t,AGQ����`_�(�x��8�]]V�����4l]֚�y����ޒ�aφZ!�\�I0�k��g.��Zƫ�"���	W�U,r>Q�v=˟��~����jv��"�Ղl������4\V�{'t����ڛ���F��b�fOp��c�G�5�ƌIq�b�(�ilO���)������r����lg�7<��W
S4�>5����������r����*g��qe��&�L-U���O�N5-SŶ��nݚF�`fPRF��c�y��!r��M�2HʢRa�yT�������+;���R��A@��l�Wؚ�����K!(�4�矼���"���ح�eYD���ҽW�j�)�(�%�IKz�n~��>�m�f�����n g-�F�ӥY۪7���	���a�x`�{���e����f�N��Hd�~�8=V���i�0�ea$<�n���Z"ﻍ��ZC8��󤏮r�n���a���0�)��;�R�!����G����KT>4\:��%!�IՎ��8�p��
�TM H��!�I}r��~�~�5�7�K����>ڻ&���F��uj╾�C��D�ٮ������@�d�����c CHI�7�P�N�"��X��i߹z�8_d��(x��ћ1��7UL�� :�aqh���Bv�|�^�s�0PN�ڳ�u�6x(�tPY�:�f�
RB؆�mi1NCA`P>����,4��h�#���Wn�	�zx\r�T�Dkg�*^Db���-D�w��En3ǯT^�iɋ���f�
����p��7z�qʏ�EM��`:�
z�R`L��w����uY��Y�;^P�Pd��j��̙��ר�h�wNm��B�?@�ڑ�
N���� �7m;n�"��M��m �a���v�{�j��%8U�L�x(k�ߖs�SZ��Bz/o0i��J&��9{���?����ub̃�IC�ҋ�č�x��7�2MP�!�9&�9�ⷕȵ�ϸ8P�c̮�ߏ����L*p��Gf�|�U�\G �8��>���Gn���ġv���%�jR0�W��M�� ���'M\�S'X	!���AJN�,}���aIX��ca�V([7�sğ��X	Ƚ?�0�T�V�Km�0�i$�{-\��B���/�j�PKH I ��!~����v�x�Ib��c뚾K�p�wo��S�+N|k�	%Ŵ�U�.f}r����{.�2�6���p�-?�W�܂�4�s�G�@ɳLݿQL0����zM��h���
^��v��M���5�g�T��'٩�8���������`�_IJnUy�\�'i���W�����U@�#��^����Ix��vg��=���*�,��'��2d��۶��mt� ��D���I��^�ĉ^_r(tTH���f0�d5{���t��ϼ,�R*�������WVӲ��͉D�����-ف]|��skR��TE�M��=��Y�����O���7Ϧ��`Nr=M+���}B�;5��a����c�u������Eף 3Q2T�i���!�%<~�1�Sȱ�'�Bm[�O�KbͶN�j��Sg{�X�9��9�L�db�l����(f��b��(��HR�P
�k�K��j09��3��wd�İ*�W۽!�aW�S�	�3%~L5C����T�1a��o�m���=)�t���ٓ�!{���=u�F��듌ɾ����(3��.d �Y�a��r���ۼ���a�]lN�H���}ڌۥHUTV�+��耉��*��-ca�)%_�?4&|���#쌍\XߨxqD�b�r>߬��;��Y���9eC!���c��xl8�{B+(�bK$�똰�gV
4��͋����P��;�F,��ƿ 7�ekp�L�p7(�f��K��5����]�mU�����E͹�Y@w1�ͧ2���[}�p���*_K��v�*��.u���\��_�Y�ynl��-9��A<�f,M��$��g�1@��(yB���Is�S���A��o�T"Q�`~v��{���`�hx����-�}7�Q���c�O�B�o�E��^��y���M����ܻ��?Is�M$Y�Iǆ�:���E����r��ɺf���ޫF��aP�� ��9��e��N����������_��Ђ��$��{[z��q�Dsxȃ�|x�Ck��N�]����tg�U�:n'����BQA���m9{{�\��Q�BGY��%�@4xt�������o�U�e��f.:�Z�ֆ�mc�^vN\��CVr7���bgzI�fXr��}���9T�|N0�)��/�퀎�i��/�f:Gz�Yb�������_��\��7�>Q�?�&���84���C`�Q��v��:��F^G��A���B�i4KY0���9*6�fV��$z?Ì��[���-����im�qY�+�������̬$P�w�1^2瑸X ��P�|�ٱ���w��W�G��v�ܥ�'�!c�;+>V��y�&;��jΊ�VC��U�>[��=b__��S5�U�0���/�0���ܡޘ��N����d�i�G�>�BH<����U|�9
a� v�i�\ഡ� E=�H�]^J�q�+�0��b�ښm�ii����<#��Ŷ��U� O�Kc[3ҟ�,�Rp�	?�J��{�����כbPA%��Y�_H�ÝoC��������s�)�o83n�C�f���*!Ѫf#�lq�=� Ͳc�_�_>��l��x5��? J��0qi��+���oD����xL� ���Sȭ���
���	yo����$�vb ��^^���^�s�Z2��73A˛��S�.�V9���L���v����z�G�9�i��E�>*l���
��3���X#��Zn�\G�#R�6`�d�v߃K�G�P��y��5��!ۊ��X3�8�A;�!cǝAY9�+��z�y&q�5�\dW rP��^t�&3��QEh�Ȧ*���x:���?�Y���^6�bb�s��A����M�����u*�)���}�B�[i��6X�$��=��D3�y�+/hn�pP:8R
b��@�	�@CgB��$��jŵ�P� ;�x"�b�p_=H<�i����_eV�^�u֣@�(�%|w�'�Q�	��<�.���S� ���L,Z�zI����l�&��?�){�I�)!2g��)�;}p��e��(�t����p�ߔ�;��ӫn@�pR��ƀ{Q}y�iu�ڈ}g"�)Y(�k�/�m��x@»���.i�Ѭ��� k$ﳵ�V*$EF��m����ӏ�j ۏ ։���4gm�K��ỵ`�W���}i]�����<�|�~��ƻ����ӷ�!�i;�%�A�y� Gu2},�����83�s� ����Kw�6��?���5!�$o��ϯO�(�Q_����*+d����K���@Mn���;f��ݡVrJ)�ŭ�4��	�,�t��~�u�	T>������D�����T`b§�����{G�ϖ��Q�=k�.i�y���S�9�bk�)ki-BF`��a�d�j3���YG}m%�5fM
$܀p뺿�/׆W9��*}$uZ𶜅ކ���Zф��B`�э5� �,o� nJ���Q�1mK���cM*���u�p�%Kmx�c�����j
=
��ۤj����쁼�?�����C7]Q�rSmNZto��1�]�}Ξ���q#��C���7&dZ������$R�?܂߹���I���,:��c��$�ADD�[L�Z:VE\h�? ܐG^ ǰ�[�O���#G���C��Zb*���E�"0�� հp����ڊ��]�t))�������;�h���N��s�@�t ���
�=��j�g2�ǣ���P������ ��eha&����'�B	Lؼ�����Z�;�㔁LSx QvЁ��*>M2h�t�l>-�zʬ<�.k�;�},�j�'�&T���=���6�D@lĖ�y�O�W�_�E�����󎡒�b�?��,^��.�~C��v;P6���W��?������.8!�/Eҷ���j���+��z�O�^��פFE<�i�*6��Q�r�T�����d9��	~�;B���-�C�]�s�a��T�G�@ҋ������:�h�r���Z�̈́N��Q���^'�'���� "4F�w���2щ^C�vыp��D#g^q�p�4h�8bk���h_P�E#�%�sK���;�8�d-Iw:�;�?�y���j���J��w��u8�@'����U����̙�S�=E�آ���d�h
u�Ә���b�PkNQqD�3-�����XB�F�q����@�9�X�Y�Ov!3��RC �S��ʯ�� 15�{t�+�@ny�l�#�mX5	G�����b�2�-*5A�4��P�u�9Z�@d����p���ݷ[��0tn�V�S��֡��a� {~t���/8uz�턞F;6��&G��(ʬ�>e>;|D�"K�)0�ć�`�O, Tf�X�M��Z���9">m�i�94�b]��i#�����h� JLb��O2b2"�����VHP�$��[+�d6���j�����Ɛ��8?B���a�kq�����ޑ�k��E��aܻ�8]gH��B����x�5m�Ԕ%$�r�ʃUa����!-N6�F�N_��2t�y΁��_��K�w�` �$p�1�9]�E�q��Y�C�z�0(Z��M���̓$�`=����y��VHM.���!J�3~2[7�ҐmJ@�Q
�ȃ������=Bճ�߽m%q@n]�Eh��]�¾�޷�)�x'�9�-1��E"�%��i(�n�6fr2�)��תo�WƝB�&/#cץf�]�s*ˮ)��|�}���3C� ���o=� ���i���e���
��ꉼ��򯗮��3��y��*6�M�@����i��-����e퐸sݗҶ�Z���w����e�;]JK���׈�N7�����-/�O"��|\[P��rܒo�j��E/�p6��K暑z�;#BD])o��.�Q3`/+m�	�o֮R[]G�qIH�|qBo
H%}�S�t���i[%��L<z@�)6�d�����~N2�I��CQX�Te�(�A�'<�� աM@1"��3���3�ʭ�	����K�	�VN�h<1l�s�!�IۦcC���-[��Z��!38 ܫ8c�ya8A����J�!��d�*�Vf�Cc1\����$�"�sV{�M�!�%�:3> AZ58�d��	�;� KbކM!�g�
W�{�T+� c�h%�i�m�Z�q��W.L\mV ��_u��(L�������]C���\�W�P>vT��������z�C��3?Èu-������]��(xU3�^Q���@$�i�ڄ�}��D
�h���B��H��M]��:��9�5X}�����Zv����#� ��ف	��ׁ�2ap�c����i@��/D��(f���s=ԅr�TPpP����?�s�*f��R3�){B�>ŔQ)A���l�̓���t#��EY�鵌w��2G�BL��# �ɗ�>2$��6�T>`�a]�n�Z}�?�D����mK�;�܇��<��dl���S{m6w�D�xd1������'����wW5ڋ3��I7%�`X�	�śU�����3�}&b�^��+���� �.�����X4)6�d���o�x�0��������&��>�ɧ���9ɧ�����۰l���R��R���=b� ���e��I
�.���9=�r�k�a�E��)�Vj��.�H�c�@����D��Ǿi(2Tk���S���L�[	���U���>��m�B�ʟ<������O������Ű�bh�R,Z|��
.Dʎ�[�V�[-^ә2W��*wchE��Zo3iɄ���t����?:��:EV5[��8�ƨk�ˤ�����.��dO��fz��0�󙘻����cE��D"w�NǙ��ɔ��g�-rշm$�jx���wz%���ڭ(mԴ(�uak޻�}���XVA����ʵ��6��/�ͶQ0S4����N��9�Ü)UcP��M���dq��S��26�q�H���K2v�;_O�0�\�D:�'y
���.�,w�po����w���D��8Km� �p�9~Cc2�/h|?�����=/�<����pK��8��ϖ��-�Sz�����3>�KU�?2��^S�e�%M ��(Ë��5J�U��J9�ٷ��]�^%ٿ�`���a����ݿU�H����>V���)
��$���^篯�Y N��0�fG����45A~�;S����rf�g����nȿ��ǭ֩^�(,1G�b'��������8WKsZq�9���t.�4#�[}�f��t���Lj"�;���f��*�a6uz}�e�9|x�I�9"Z�P�;�J��\R]<���Ol���y\����s���;���|�Cq�e�fdl!������,[��}�$�)=zӋ{[�Yr�'6���Xuޣ�Y�n�t�š9&NioɄ�72�r������%���͆-��U�7c�,���屃?T�JE�
Sq�E^��u��(�d��ͻ;��F�P���@7�X�0am�����#.0��%Ss�%5���^$�[1k�"[&�O��e�`U�����b�m_�*F�9A䨧*$1��BB佨��|M��zq'R�]&�e���~�-s����[� _�t�|�gz�2�0��l�T1�E0o��H���R���F����T������QF���d�f>:�)Bh�_�V� ��
�"ѩ���2:ܘ2x#��T�ica˼�����I6T��2\qݪ����v/$�ɘ�iܱ���ѐ�c���9��p�����*⸥{�U�����"N�j�N� *��ߨWs����&�G|�l�x�;�P)y�j���0�DҊ;�zvy�K����Ǣn�lo���
��X�G֨ܘ�{6�o��Q#���O���pv �n�H@5�vh
�U�����e����u�@y�+I2�<l�oG¸����7 �5y�����+������@���� �ܧ�h�?�DH�d	�L,d�:'Ka�U����A��2�`5���Q�p�#�6ےz)md�f�H�Oq%��k��B	3i"�Ȁ�ދw����Fs�0��3R��b�;J�9���E��>|�3�C�k9p@�Z#�eYWŔ���\C�G@Cwf��_Ob�O7c��q�+��a�\��L�g�Qc��~�)�Y�����NEW��u�f�z�2�X�ũ�J�oD� Z�P���׶<���Uf�����|M�heC�A����|KJ��t@N|�즅�<�s:�e/�7p��J!�,���^�'�:P�vVQ3-��3z��^<7���>�.E����"T>V!֤��d`����.��;��k�;5��"��Īyw�� o���MA=
̵
]qW�8�ݟ{S��X�@b8ۥt:�b�f�ܨ�x�LG��t* ��B���u�Ll^��v�;[{I�`�ߛ4�3	̕a����X/6�7r�=��jV:FQ>?-T�Λ?6���~�c���*����,4-;k�	FY���Lڦ��j����V�"[M��,k�]�!�Ѡ]���n=���Er�5��,�3�������ɍ"b�տ���/�w1����g�'r#���[hr%g4�\����g�AJϐ}�ZR�x�q�w�z>�Q�ӹ`�ń�F�n�t�#cJF�Ȯ94o��i�c��m~�ֻ����:�.5Z$ x�k���ݧ) ����Ji^t�hR����Q��Š_��r�w���3�LWk�K�ؽ��������L;�-xT���p�]��ƨ��n�jAZ��Uo�d/�b��ܡJC���l��-��q�)@���/�5N.���:&.(�'��m�pv27��y�"DN�p햼���#!p�%�P^s͵�$f_�*C�Κ�*���;�(����URHwU��J�ˊ�C����	L��,��htQ�d�_�#�F�؁)!��-]h�oGU�����.�H��V�t�r-�~e�F�\b���H+����Ƅ��//�OŠ���
I���Z&� 	Mi<5[;�"xV5�I{�m�Y���4x��.�1�����I��s��p�k�8��Ht�@��Q�_o�nA��mn��˴Æ����l��!(L�S(9��mJ�Ⴗܶ��c�	f'��?�2����Ƹ��p��<�-���e�)�Z��Dpy�OXf=<;Q�@��|*�c`铋��Tj���`��]��f�T
�~)�a�1 �-]๥�>>�b�Q�/����e���'�����|�Qgg��2��O�`r���Z��i|��u�P7T[�B��J��DP�`�>�֟p�
�vO���%mWY1�-f)R�9G�IɌ��'?��ٍ^�e/���G	����J��~ ��m����Ŗ���d
ԿH�AT�n �vܹV�B����+"銐��_*�9��ɀ�AKzJ l�w'��Cnz�����޸��:�e��L<�~#�bV�[����dO�P#���F���|
�)m����7֖e�y����.u�Þ��`�ɣ�����p�b4[�z��-)D��Cw���o"�=�M�yF#� �nSxE/�^VJ5��?�S@?�%x��������2�<x�8XW�������̕dn��,l��Y�]�r�+L��������8��&��r;C��7'� �z�������
����(�T}�%���&���8
�d�t G@���&���8X"k�#��hk���2��)�b�HO�Wh�A�의�9����Þ�		�ҩ8�m�-�]֐-�ovPze��4�\6ƥ�8��Ym´����KP����m���k�"�x�O�*�ZAr�Ll��]�$��� ��m%�}]�Ae�(�Ɖk����M�M6,^�Ŝ��7�|�dhK?CN��~b��#r���XH;��H���]�}hG)�ӌ#��9�D-�)z!O_T>�����¨�4��2C�����b;^����	S�X�1�x,Ë1�jYi>g�Rn���dߨaITq�B��Y�?�Hyb0�����=�ܨ��az�W�u��}���b�fCo?·���� ��sZ��(K���V���}1��GסN&h(LxT���ƴMp�K,V[|ƫB�^�G0L �p޷�@��A�����fYq���Nҕ��nY����(�oE�)�DoK�D�?�:���*ej}��N��:ۧD�	�N$�E�i�O}�4���f�J��@����}���MR��Z�Zy�K�
\I`�������n�yRA��P�GR�{!���6M	$�&2a�����!{�g*�s$��4'[��н_6�%����Ճ�(Y!�c��@^qNNE__um�ލ��Ʌ����1��_�����Q���I<NM�Z�	Ge���F���-�@ �v�Cfe�6�P��~��t��+�:��h��WBi�!l�����rqR5,�ԩċ�{��=�BMQ�¹�(�R��h��
�]r
k�D�����r&�t������i(��Eۀ� )c��գ�S�'�{8EHvn�>;����Mѯ��QICzOzZ�e6��^(�{{y8q�Hxj��;�������8/Z��?��M��.|x���/��
�����F��g3�{����U��Xzȁ�}~�GD;[�5����EO��u��Vc��"�6��YY��	%�/���i�y4��@S-���M��6�Ym-b3b	W�����h���-ߓ����A�eW紣��{'cA��8�m��ۜ�Akɍ��yw6���q�K�kG��W��4�\΄�d@�d]�.��ƕ� �8#���ؒ�� ���\3	N��\�t10�}�Ѱ~�C�?7�k���pTJ�"�#Ѝ/�[ŰUk6B��BO'j����3���k��\�8<K��5*�C'5���9�Ӊ�b��K"(��N�d�/:����b Z�߆��]�xP)J�%��EA��
1�Tu�<�.��
� W��Bu
O^`�\�p(�>���.�[��>�]�4��[�B�D,�0SԒC�1N�J~+!�rQ%W�Wx�t��� �U���l[9�����M昚�������;�S�.��.��E����Tm��`},�	��`l}���[3�Ќj��tL"dy�X��@�ewj=%�k�%,��r�TW��(f^rn�R����L{�b`�6;e���D��a�Y��z+s�Gm����-�(9φ�3j@��_���#�P�P�u��w����j�� �N��uhDJK�,��ߍ牰3�h��/�\sit_c:n;�k�.��Gy���y��g)D���f�"�3�!�DQ!�t�o�[+��1���]�(�9Qcx{�+��C�6�S���f�r�mb#-����>c�K2��v����L���ĵ�ͤ J�lgv{�W�T�]`���-���F=�Gyl&���QM?�j�H6a%�Mk7Tи{��������D�!$�8�e�5+���o��������T�O�GE�3�&�H�F���pyu���<��A�0O��l3��{ZZ穟Z6�Ň��WU5"��-0�-\A�Ќ: s�!���l5Kf�"f��N��D����A�EA�b�����J�.I	������un�+����p#�66b�A߶��t0�.�t��T���E��ﻍ3*�!օ�x��EZ��ҜB���#�ǽ�j��:M�}9��%w����{�P2P��+a���\{l�F
�"%���at��m�w�t�5�^
y 4�k��R������B�Ϋ��^P����;�t�;,I�L��;�@auO�jR�L$�º5�J��1�a���о�::���+��&$g纘L�*�E��B��8��!n����ՂiǙ��H������]���ZܻD�Y�j�HDH`��?���֯A��X�%�����}?��i�d�q^�F�/�
�~U���
�ޖ3,U��{�����;��UhN%���3� "<�w��O�5��S��&�h�0\P�͇v�=^�K6c��!��*b9�&",58xῨ'x�/y� �1��c�E��g���㰽8 �:W��X$�:���ȌQ܌\���ԲN63]0I�o�S�S�)���y�P��1�) 2��fߠ!�-����v���Rz=b���D�T�ٖ_��j��<�!B=OܥC���!I� �R.*�/^+;M���T̺��
]z�yK��y����`�T��-���bKMc��< ��v2)�x+�q�0���s�ŀ�b,"�:z��oۃ�����@H�|�&��*����∪�8�|Ax6�7sP)ls4_��XB�UВ�{�r��(p�]B����X�A��l��D3���3��?OOz=K�U�P�N��
5��	$��˗e�T�í~%.��[]�3���Ax�#��*U��yC��+P���mi�ƃ��h�x̎^70q��I���T��9H1v��=�h���l����o��SҞ�4�l�+�ǁ��������M_�E- ��<	��۠���L��]�UFJK3�HJH^�P�'�[��%�Q�]4�-���}�歷��ƻ�ah�u�H�F�D�1���� ��#w�SZ�	����C��e�  Pe����Q�l�/x��iM������ʬC��ud�I�]`�x�#�&�;&��8��L_�8����Q�j�Uf1i�Ip('|�  �fd�5���7���9#[q�"�O�(��c@��c�jJѓ���ݖ��'>���xl�9��oF�w)�IM
�˹o���?�H�"�A���M�a#�7D�/E^a4K,N��oH2�iE��o�9�
;�VzT���Ll�����{�Si��;I�.��V�_"*4��b|����{�l^���VD�6`a��y����p���#O��|{w��o4R<���T��e��p��}�G^^�ͪ����*��d��;�|.?"�Ӹ!=d�%�{��ã�|u�hCy���������p+�o�ީ��E6s��TF+ܓ��)i�,ǒh��|��c����>� ����9�=���FŪ��c�w�h�7�r����i�@a2?�IJĭa�V����V�~G��{f�=5�xm�6@g�/����!���m���#2�(1n�x�6����$He#\F��J���wqV��n��������v�=#����
���λvt�u#��SŦ�>J��&�"�G~"�OĂ�d�R���e,��#[�l(�x��'�D*��Ӱ���)��Z��|�CԛW�91'��V�|�ҁe�	n�G>���^:�����OVM�a���|��gL��gX����I�(['�����J�_�1��LBPɟ��z��s̈�2Y�	7���?$k��ם1BDL\��כz�N&���]o���\�\��zmd�����;���(U�:��q�#�@�
���/l�2%w��1����!���f"����l(�L���kX�� �%EW<Yl�q_R�
�:���?�<`X�]�ѷ|��o=s�B�+��8�י1�V�a^��̤��yMH�ذ���HH�;�[�)��a��Dwzd����E�>�� ���w��� �qw��z��<
Dg���c�.KQL��$RE�uS��У��5��%֨��LU����#�W[{2UH��,���VLoD�:[۬�xYF4 � ��������V����&3�YJ{��C�Y�I�	��!��W�ڨM)�NB��ϕ�Ċ���y�Bm��t齖^p-{��e��j�7@�j4f��JӇ|k;
_(Z�q����O� >�/&�����Si��i6���<1lEd\�\r�.``��̓��&!wګ5M�LA>K�tJ��Z,c�������'Q����"t@Z�/���f��z.��"�2o�Q�Mϱ�"��k�ه�����4�e����2Փ��Q7�-���̑^{7Q����y�����V��ڛ���0*@��D�X�[Yms3u)���;�2>g�yk{DtK�%h�.�p.����g�D���c�S#�Kv=(���^ł-%��wveЕ���$d��7d��Z8�R�a����l��$b�l�.ف��j�*&�xM�aS;�H�r��uv����q<���M 	�)7�U>���fiXJ(�V�iq�<o�� ���a�:�z��Ӹ����O
"��|F���H���v��Z�|�f��i��&Gu+�l�>�[�ۋ�l��۠|�ۛ^���>�-{a����c��L�����E���Jrs�qS��s�R�&]�-&���Yz���L+'�eYj�����r&���1��!n-k�?�hޟ�k����q�jfss��V�Oؑ��-�{'��UF_H�fA>���:�iL �d�b�s?R���I���'����.\6��#�f,�[�g�,��ft���kӛp�Du��A����;t�dژ�'k���S�կ\`�J��(���M�?��={�XC?���S��1�4��
inN7(b�HGBZ�g�pҋ�.���o�S�w���ێ�k�-3mKWyPS R���d��8d�Y2?
�e96�L�Q��IL}/:��kk�R=��Ox�N`�z3�d/pY喕����#�813<��P��(sl��I�(
<8wW��ͮ�=��
hxjrJѽS�?�%��A&ǱwT��w0�\V�&[Z�M��J�C�h�^�����0f7����S����Es�:05|�К�g��(<څ}L��N�q1�����?�/$��ꋁ��O��۬zdO�/�,q2A5G_E�ΝV�y��{�����y�B��{�4R�La��WA/�����Q�W���)�
�N��Y1�h�.��͛�����C��D�$�p���(�wN���X}.ah�ժ�>�	����<�ȈL)>|��F�����@�:K�R�
�+�C5����g�p7|��sCc�f+�Z���*�B���W�A����'S�v��"���qJHw��>��8 Sҡ�ʟ\�_.7���s�JDZ��Å�8u������cض$%�N�j��H׬�Lep���d�5o�"�&��gul�Ob������#P����l���@��4����̌���f��U�i���������0���)op�dŧ	V�D%)~�.��:R���b�-E+��,S}x$���[ D.�j|q�e�,*>��1�>��C�P[�n��^�&�ǫX��"�n�dg�H�B���6���ξ��b|*`��x�*�w�pZf[��"��zb
�SoU�D���b�HX%��G�wS�6,`RT��U1��G0pZ�x��!�{�W� �2��xl��ݘ�d|���Ɨ���#�9���ͅ@�1(����|V��A���{8`	ٍ����ϓH�ʓa֫����nĩ+�)�t~7�gG���)��m�Nԣ��~?����}�����cW-��
�d[��#�ye2VIa�$)����6������~�!�tM�!�R�143�	���	g���_m�Ra�6�H�~f���g?���A]!UJv�mi���3����8�a���8��d[
e��M��ZN:TS��tr��|�_]@́�����h�7Z� {d\m�N_�} (��z�E@���hTE�p�/��m`AX_��qHT��� ����\p��)�e̒�WW�x����li������]ɐ���d.�OӴbL%�ؗa�`��)@�"�B�E阀F� �c�81$� ��~Y����p�������M�Ħ,������<��r.c��=���ʔ�����v?0)�kRav������)q��:$L0�6���*x����y)��DP:�T?n�eL�HM�4~�)�$�m�q�PlwE5�]D�c�(h��/��u1�K���n� ��J3b�����cu��c5L�A�����.%��M5K^�X��K��%rݾ�Z��Բ�&�E��A�wȢg^�h���C�jѲZ��O��8�����i�ؔ"��ê�	�4�]�Y�/q3��{$V���?r���1e��CF�⒝`>�@	�a�{�s9�|��)�3�-dٰ%�	�`�j�2����̺Ov?���|�[����ʁga��+s�1V�B��akt#树���a�,� L�ЉNy������6>c�G�*�G�Ҟ"�I�BW�x���}k����)�L��©ؽ�T���1U�$$|��YiV��yS��nў��Y͸金��dʚ�#2L_��$�0d���5t�[Pe�eS4j�f�>*7Z��k��!�����(�B6~u�	��u�L�vÿ B�D\�RID��<������
d��=�[D�cO�gďpܢ"k�^#�-�]�q�U� ��z�7�[���Bf����2p�u�>[o.�e���e�$�%�������0���k�{���N�k����~C�~�Z�:6Wc�:%�\`�j�����m2�y��� ���Ga7�?8`�w�����z�&��dTK?6���J�[�i- e/~<K0�����W��T-��[<sj|%��;�����׻������-l,Ҋi
2�9���+HH6�k��a�kK0�Dp���c�O���x���u�b��l��RF�`?X��d���}Ǉ�'p��ӶY�ࣞD{Z���v��O�����2:�ox���=���os�l�L����E�gU��ZY`�<�����rن���3��,�8Vdr�2Or���8�p~�����u��A���:�n�����?���V~|�#�cߓ}�ůa�u#[�zh)peo�`r�ώ�ѹ���;4m�]��_�5�Y0s�k�f������2�ݷ����LY�\�w�!�j�ZCTҵ��JڤM\�I�e>���t���/��ċW!xB��؟%4u���gZO �i����W(�ܶ��pU�K/�����
�HJ{)��Tf�~K��~�4�f*���}�q��� ���@�|el���!B�+���/�g^���<��%UY�Ǡ1+�8"+Ь������蟝� p�*Ǻ=��к�	�T��Uz^�������<�6�"j?U!ă���]�)�n�P.��Y�4i5;7mF��X������T);��Բs)�&P	���'�\%�r@,^M�,Ee��I*�rF�5���Y�ӽ���3X2f�=���-�X�(��� .+ݭ��^�Gjڟ0 ubb^��s��ma� ��X���pY��C1QʼN|���!���vdrB^�1��f�2ԅp|�!�+MH��B������&RTӮ�>`�E��u�J�=��6��Lڻ}�D�����g����ߎ��>Lr���4r����ي����V�G��
ZLe9�u�t��L?�Ľ��s������Xk��0oUܣM���'!ؼ�b�R�vֿ�V�������q,������YWT�gt��/O��gE���D����_�u�,y�xhh�� Tw�%�r�*��2�����И�ViS�֥ԙ$�on����X��Cb��蚩�A�����>���Dz�1��y�R�J>�+����Lށb��6�O�_�)�s�%DG� j��M����J����#˜�<������h�_f�>+7q�,���a���:+��C;���}�b4����g�����Y���X��Q��Ɇ���A���运0�{��,����T܉���YU��&`9ա�c��w�mk�ǈ^����2F�����K�����ϸ~����o����͊V�8�p������x�������%�<)]|\�KRE ���z��pt�=Z-�<
#�J�S�$�".�w�%�,��v�m�B�iH:���\2�4Us���i2|���2�F>�|�h5F˴}y�����Q��C��i-D�9*}HIљ�R���u�7�a�����,)A��"bu"�zhf�� ��қ�y#����N�xh�b�n�����ܓ����߻�d_�
}W�����ס��%�&�yS���(Z��:j�>�����P��*~wgL}gQ�֑�El}3#O�';"]�UYY��H4��Ճ�-�b�g�~f�ep��i�����OT��/�+��s�/G�Y��:�hԧ0n��{ͤO�N����:*;qG3m!���Ļs�?�f"�J�z��Lbs�[��&�:"����|���]����
�g����<_�n	7(J�4a<�#��XFi�lǪ0��:�EJ�դ	gיQ�S�o����/� �w9���i��\�R��i�(2��)���n�Յ,6�יc18�K Kl�<�Vx7�$��$$0 ֬C�E���J���{|!��j���g�|�:��8E��e�/�]��z,Џ=�� ȿRW���ס1�g��ީ��f�m�T�����)D��J�L��] >��^�t5n�~9Q�R�� y�v;�A��9��anR鬂�[�4`y�A�ۆ".���U{2�}�D���[��ҡ�-)��8��=��%gQ�M��`�A���	��.�~1���F� ~��a>�Qˀ��Fl8�5jN
4���})2�(�ۃ�A㜁w��649����Լ��x�\Y��R
��F�]ۄT��V��S��vO�"4�ǿ/,S����������e�=aU*���?����;�/xW���ˉ��L��� ;��}z�v���&Q"'����w;6M�z8a��K8��U�}m������+i��Rڭu26�n�?_�\#)@u$굦�����Gfu�LzI�v2�cj�5��9HB����֋v��ΥG$|����^#��.���w�s�K���ا�q��)��������b0'�:�#�S�1j�X�(Qh8�՞0�֙!�f��ߩb��K�4V�d�Cs@ˋr�}N�|���Ҿ�`��Daa��fttwJ<�U5���hPy�b|:��~�r#�L�=e*O �-��Z9âӥ ��94����0l��6��YE��,͒k�Y�<�,[�8�(�2QJ�' ���+uʡ
�D�P�)հ����	�jB�,����?�����-����:�����!���m T�2;�Ό�݉���*SBA���h(D��	3�}���H���Ig�X ����	�Fq���>4��a],����Q]x�N�h�AX��	fٳ8*��P��s3�p(�j[W+���M��D�(c869��!d`��}�m`��\���x���O.��_
�m�e�V�hx<�Z.�>\�������}����I�d#�_R�f�cGAU�� 7w���\�𭠑���2�����|��wq/���q�4(�� #u��wu^�'+^�Jr}�@���S'�S����f�( 5#���w����p��=�C�g:1�nUӾbM�	����B�,3BW�59K���
췦�ԡ��@G����8Fl�`�������x� �-��ȧ����>�q�v%�n[�{�ҝ@�Z+�嗌30�Us�'��S�4��@2J���"_�v�S��TW�ϺY�������7o^��E@���cK�������)��7pF+��L�xټ�	,ǟ�ǎ/#�wrQ�FB��=YB�n��|�?3�f�;�?�p��`Q$�u�[k�����^t��ņ�My>4UPR}���cy̛ؽ�<���2 �y��6C����8f(��F:-7F�?�)Ƚ�6�n���,�g���6E^nV0D,�V��b�O�e�Z�AM�n���[��-��L*�@�W xң6�Ʃ�/<�6F��e1�{@0�l����*���� �\� ��T߈u��C��Pu���+]�6A�՜�oCo!�+E��G����9X�cC�xKZa�12�UZ+�H�W�2��	8����|��%+ y�?��~m�<���o����Q��X�
Ti��_�����Z�^9��#��%}3h���A�$����=���j2�W�v�w����3A��4BZ�����Ǵ��a�h���s1}��<@<X��(/y����dbp��Dt�!ȍ��;�h
��]��w@�|#ooS:���0OZ�(K���'ㆃ	�4�%j�x��]d�k%*�U�8(����e�,����c�d�Z�(G��6>P� �`��m[7�lQ����h�l��r�uE�R��C�I��E��lm7�D�0�\dGe>8w
*4X;0�S���PL����B�f�C8\^��_G�:\7��Yt��7�0M��~J- �(̍��ʋ��q��B~y%�b�=���U�j�́B��D�K�v�^@	�RuHB���:G�� UB'�U~EQI���r��Z�?'d�ޒ&ꖶ[@���R	Ȟ D�{�t%�SL�T%Z2�&ս��L�8��/e��1���J�8�iyfa�o6
ɼ,�iN�4�ҳ�:��8�dU��oyo6I�.�������%� aK,H�$��k��nHL�~_S	6�e,�E�~�!i-8���5�YY'���(���tT���O�%�J�%:�K��8��,��p �Ҽ���-X��gF���_T�=�b<1q�#u���sy9�� Wj�:6��1����N�\0�YG�t!1x.��^� ���/��F@�h����U���&a�v���9ߣ�
���'��o6��FI��\!Q���=#�p�T1���s��bv��f��EC���8�Jwfft�� r�!�e��C�$�4�C9��;��ˈ��� �1_��
&L�o�^���_�����Q���Hb�>f=&6�խ��
��X�\2�pO��E处�=(�/t�c�j�겊������./,�lؠ4���aE�6V��17���)7.G��fMk��0˱��.��������.Y|ȍp�=�T,V�-aT"�Bs�|����F��Ɨ2�_��ȾE�v�2�z��b��0����G[���Z>w_��DlY䚸���N�^��.�98h*J�b�E&��<��~X��� d�7�(��3��A�?�T�`���iL"�}��f�s��-�_9��O�����݅��m�M��2��hS+���/���.2|E��zeD����8A�~����&WF! p���}5��5u�k�7wM����,�a�R��p��ƊȀ4��Ҋ�Aغ���mC�-�7�1��� 5��l\	+2,
���bdB5